/* Automatically generated palette ROM */

module palette_rom(
    input  logic [7:0] addr,
    output logic [11:0] data
);

    parameter ADDR_WIDTH = 8;
    parameter DATA_WIDTH = 12;
    // ROM definition
     parameter [0:194-1][DATA_WIDTH-1:0] PALETTE_ROM = {
        12'b110011011111, // Index 0
        12'b000000000000, // Index 1
        12'b101110000101, // Index 2
        12'b111010111000, // Index 3
        12'b100101100100, // Index 4
        12'b110010010111, // Index 5
        12'b011101010011, // Index 6
        12'b101010000110, // Index 7
        12'b010100110010, // Index 8
        12'b100001100101, // Index 9
        12'b100010001000, // Index 10
        12'b101110111011, // Index 11
        12'b011001100110, // Index 12
        12'b100110011001, // Index 13
        12'b011101010100, // Index 14
        12'b101010000111, // Index 15
        12'b011110110100, // Index 16
        12'b101011100111, // Index 17
        12'b011010100011, // Index 18
        12'b100111010110, // Index 19
        12'b011010100100, // Index 20
        12'b100111010111, // Index 21
        12'b010110010011, // Index 22
        12'b100011000110, // Index 23
        12'b011110110101, // Index 24
        12'b101011101000, // Index 25
        12'b010110010010, // Index 26
        12'b100011000101, // Index 27
        12'b100010110101, // Index 28
        12'b101111101000, // Index 29
        12'b100111000110, // Index 30
        12'b110011111001, // Index 31
        12'b100110110110, // Index 32
        12'b110011101001, // Index 33
        12'b011010010011, // Index 34
        12'b100111000110, // Index 35
        12'b100011000100, // Index 36
        12'b101111110111, // Index 37
        12'b010110000011, // Index 38
        12'b100010110110, // Index 39
        12'b010001110010, // Index 40
        12'b011110100101, // Index 41
        12'b010101110011, // Index 42
        12'b100010100110, // Index 43
        12'b010001110011, // Index 44
        12'b011110100110, // Index 45
        12'b011110100100, // Index 46
        12'b101011010111, // Index 47
        12'b011111000100, // Index 48
        12'b101011110111, // Index 49
        12'b010000110010, // Index 50
        12'b011101100101, // Index 51
        12'b100101110100, // Index 52
        12'b110010100111, // Index 53
        12'b001100100001, // Index 54
        12'b011001010100, // Index 55
        12'b010101000010, // Index 56
        12'b100001110101, // Index 57
        12'b101110010101, // Index 58
        12'b111011001000, // Index 59
        12'b101010000101, // Index 60
        12'b110110111000, // Index 61
        12'b110010010110, // Index 62
        12'b111111001001, // Index 63
        12'b011101100011, // Index 64
        12'b101010010110, // Index 65
        12'b100110000100, // Index 66
        12'b110010110111, // Index 67
        12'b011001010010, // Index 68
        12'b100110000101, // Index 69
        12'b010101100010, // Index 70
        12'b100010010101, // Index 71
        12'b000000000000, // Index 72
        12'b001100110011, // Index 73
        12'b001101000010, // Index 74
        12'b011001110101, // Index 75
        12'b011010000011, // Index 76
        12'b100110110110, // Index 77
        12'b011110010010, // Index 78
        12'b101011000101, // Index 79
        12'b101101101100, // Index 80
        12'b111010011111, // Index 81
        12'b110101111110, // Index 82
        12'b111110101111, // Index 83
        12'b100101011000, // Index 84
        12'b110010001011, // Index 85
        12'b001000100010, // Index 86
        12'b010101010101, // Index 87
        12'b100101010100, // Index 88
        12'b110010000111, // Index 89
        12'b010000100001, // Index 90
        12'b011101010100, // Index 91
        12'b011101110111, // Index 92
        12'b101010101010, // Index 93
        12'b001100100010, // Index 94
        12'b011001010101, // Index 95
        12'b000100010001, // Index 96
        12'b010001000100, // Index 97
        12'b101010101010, // Index 98
        12'b110111011101, // Index 99
        12'b010101010101, // Index 100
        12'b100010001000, // Index 101
        12'b101110111011, // Index 102
        12'b111011101110, // Index 103
        12'b000100010000, // Index 104
        12'b010001000011, // Index 105
        12'b011100110010, // Index 106
        12'b101001100101, // Index 107
        12'b010000100000, // Index 108
        12'b011101010011, // Index 109
        12'b001000010000, // Index 110
        12'b010101000011, // Index 111
        12'b111111111111, // Index 112
        12'b111111111111, // Index 113
        12'b110111011101, // Index 114
        12'b111111111111, // Index 115
        12'b000100000000, // Index 116
        12'b010000110011, // Index 117
        12'b001000100001, // Index 118
        12'b010101010100, // Index 119
        12'b101110010110, // Index 120
        12'b111011001001, // Index 121
        12'b100101010011, // Index 122
        12'b110010000110, // Index 123
        12'b101001100011, // Index 124
        12'b110110010110, // Index 125
        12'b110111001100, // Index 126
        12'b111111111111, // Index 127
        12'b110011001100, // Index 128
        12'b111111111111, // Index 129
        12'b111011101110, // Index 130
        12'b111111111111, // Index 131
        12'b111111000010, // Index 132
        12'b111111110101, // Index 133
        12'b111110110010, // Index 134
        12'b111111100101, // Index 135
        12'b110110010011, // Index 136
        12'b111111000110, // Index 137
        12'b111111111001, // Index 138
        12'b111111111100, // Index 139
        12'b111111111011, // Index 140
        12'b111111111110, // Index 141
        12'b111111100100, // Index 142
        12'b111111110111, // Index 143
        12'b111111010011, // Index 144
        12'b111111110110, // Index 145
        12'b110010000010, // Index 146
        12'b111110110101, // Index 147
        12'b111000100000, // Index 148
        12'b111101010011, // Index 149
        12'b101100100000, // Index 150
        12'b111001010011, // Index 151
        12'b101000010000, // Index 152
        12'b110101000011, // Index 153
        12'b011100000000, // Index 154
        12'b101000110011, // Index 155
        12'b100100010000, // Index 156
        12'b110001000011, // Index 157
        12'b010011101110, // Index 158
        12'b011111111111, // Index 159
        12'b001111101110, // Index 160
        12'b011011111111, // Index 161
        12'b000111001100, // Index 162
        12'b010011111111, // Index 163
        12'b110111111111, // Index 164
        12'b111111111111, // Index 165
        12'b100111111110, // Index 166
        12'b110011111111, // Index 167
        12'b011011111110, // Index 168
        12'b100111111111, // Index 169
        12'b011111111111, // Index 170
        12'b101011111111, // Index 171
        12'b000010111011, // Index 172
        12'b001111101110, // Index 173
        12'b010101000100, // Index 174
        12'b100001110111, // Index 175
        12'b001100110011, // Index 176
        12'b011001100110, // Index 177
        12'b100110011001, // Index 178
        12'b110011001100, // Index 179
        12'b011001001001, // Index 180
        12'b100101111100, // Index 181
        12'b011101011011, // Index 182
        12'b101010001110, // Index 183
        12'b100001101100, // Index 184
        12'b101110011111, // Index 185
        12'b110010011111, // Index 186
        12'b111111001111, // Index 187
        12'b111111001110, // Index 188
        12'b111111111111, // Index 189
        12'b101001111111, // Index 190
        12'b110110101111, // Index 191
        12'b010100111001, // Index 192
        12'b100001101100, // Index 193
    };

    assign data = PALETTE_ROM[addr];

endmodule