module cos_rom (
    input logic [8:0] angle, // Input angle from 0 to 359
    output int cos_value // Output cos value * 2^16
);

    always_comb begin
        case (angle)
            9'd0: cos_value = 65536;
            9'd1: cos_value = 65526;
            9'd2: cos_value = 65496;
            9'd3: cos_value = 65446;
            9'd4: cos_value = 65376;
            9'd5: cos_value = 65286;
            9'd6: cos_value = 65176;
            9'd7: cos_value = 65047;
            9'd8: cos_value = 64898;
            9'd9: cos_value = 64729;
            9'd10: cos_value = 64540;
            9'd11: cos_value = 64331;
            9'd12: cos_value = 64103;
            9'd13: cos_value = 63856;
            9'd14: cos_value = 63589;
            9'd15: cos_value = 63302;
            9'd16: cos_value = 62997;
            9'd17: cos_value = 62672;
            9'd18: cos_value = 62328;
            9'd19: cos_value = 61965;
            9'd20: cos_value = 61583;
            9'd21: cos_value = 61183;
            9'd22: cos_value = 60763;
            9'd23: cos_value = 60326;
            9'd24: cos_value = 59870;
            9'd25: cos_value = 59395;
            9'd26: cos_value = 58903;
            9'd27: cos_value = 58393;
            9'd28: cos_value = 57864;
            9'd29: cos_value = 57319;
            9'd30: cos_value = 56755;
            9'd31: cos_value = 56175;
            9'd32: cos_value = 55577;
            9'd33: cos_value = 54963;
            9'd34: cos_value = 54331;
            9'd35: cos_value = 53683;
            9'd36: cos_value = 53019;
            9'd37: cos_value = 52339;
            9'd38: cos_value = 51643;
            9'd39: cos_value = 50931;
            9'd40: cos_value = 50203;
            9'd41: cos_value = 49460;
            9'd42: cos_value = 48702;
            9'd43: cos_value = 47929;
            9'd44: cos_value = 47142;
            9'd45: cos_value = 46340;
            9'd46: cos_value = 45525;
            9'd47: cos_value = 44695;
            9'd48: cos_value = 43852;
            9'd49: cos_value = 42995;
            9'd50: cos_value = 42125;
            9'd51: cos_value = 41243;
            9'd52: cos_value = 40347;
            9'd53: cos_value = 39440;
            9'd54: cos_value = 38521;
            9'd55: cos_value = 37589;
            9'd56: cos_value = 36647;
            9'd57: cos_value = 35693;
            9'd58: cos_value = 34728;
            9'd59: cos_value = 33753;
            9'd60: cos_value = 32768;
            9'd61: cos_value = 31772;
            9'd62: cos_value = 30767;
            9'd63: cos_value = 29752;
            9'd64: cos_value = 28729;
            9'd65: cos_value = 27696;
            9'd66: cos_value = 26655;
            9'd67: cos_value = 25606;
            9'd68: cos_value = 24550;
            9'd69: cos_value = 23486;
            9'd70: cos_value = 22414;
            9'd71: cos_value = 21336;
            9'd72: cos_value = 20251;
            9'd73: cos_value = 19160;
            9'd74: cos_value = 18064;
            9'd75: cos_value = 16961;
            9'd76: cos_value = 15854;
            9'd77: cos_value = 14742;
            9'd78: cos_value = 13625;
            9'd79: cos_value = 12504;
            9'd80: cos_value = 11380;
            9'd81: cos_value = 10252;
            9'd82: cos_value = 9120;
            9'd83: cos_value = 7986;
            9'd84: cos_value = 6850;
            9'd85: cos_value = 5711;
            9'd86: cos_value = 4571;
            9'd87: cos_value = 3429;
            9'd88: cos_value = 2287;
            9'd89: cos_value = 1143;
            9'd90: cos_value = 0;
            9'd91: cos_value = -1143;
            9'd92: cos_value = -2287;
            9'd93: cos_value = -3429;
            9'd94: cos_value = -4571;
            9'd95: cos_value = -5711;
            9'd96: cos_value = -6850;
            9'd97: cos_value = -7986;
            9'd98: cos_value = -9120;
            9'd99: cos_value = -10252;
            9'd100: cos_value = -11380;
            9'd101: cos_value = -12504;
            9'd102: cos_value = -13625;
            9'd103: cos_value = -14742;
            9'd104: cos_value = -15854;
            9'd105: cos_value = -16961;
            9'd106: cos_value = -18064;
            9'd107: cos_value = -19160;
            9'd108: cos_value = -20251;
            9'd109: cos_value = -21336;
            9'd110: cos_value = -22414;
            9'd111: cos_value = -23486;
            9'd112: cos_value = -24550;
            9'd113: cos_value = -25606;
            9'd114: cos_value = -26655;
            9'd115: cos_value = -27696;
            9'd116: cos_value = -28729;
            9'd117: cos_value = -29752;
            9'd118: cos_value = -30767;
            9'd119: cos_value = -31772;
            9'd120: cos_value = -32767;
            9'd121: cos_value = -33753;
            9'd122: cos_value = -34728;
            9'd123: cos_value = -35693;
            9'd124: cos_value = -36647;
            9'd125: cos_value = -37589;
            9'd126: cos_value = -38521;
            9'd127: cos_value = -39440;
            9'd128: cos_value = -40347;
            9'd129: cos_value = -41243;
            9'd130: cos_value = -42125;
            9'd131: cos_value = -42995;
            9'd132: cos_value = -43852;
            9'd133: cos_value = -44695;
            9'd134: cos_value = -45525;
            9'd135: cos_value = -46340;
            9'd136: cos_value = -47142;
            9'd137: cos_value = -47929;
            9'd138: cos_value = -48702;
            9'd139: cos_value = -49460;
            9'd140: cos_value = -50203;
            9'd141: cos_value = -50931;
            9'd142: cos_value = -51643;
            9'd143: cos_value = -52339;
            9'd144: cos_value = -53019;
            9'd145: cos_value = -53683;
            9'd146: cos_value = -54331;
            9'd147: cos_value = -54963;
            9'd148: cos_value = -55577;
            9'd149: cos_value = -56175;
            9'd150: cos_value = -56755;
            9'd151: cos_value = -57319;
            9'd152: cos_value = -57864;
            9'd153: cos_value = -58393;
            9'd154: cos_value = -58903;
            9'd155: cos_value = -59395;
            9'd156: cos_value = -59870;
            9'd157: cos_value = -60326;
            9'd158: cos_value = -60763;
            9'd159: cos_value = -61183;
            9'd160: cos_value = -61583;
            9'd161: cos_value = -61965;
            9'd162: cos_value = -62328;
            9'd163: cos_value = -62672;
            9'd164: cos_value = -62997;
            9'd165: cos_value = -63302;
            9'd166: cos_value = -63589;
            9'd167: cos_value = -63856;
            9'd168: cos_value = -64103;
            9'd169: cos_value = -64331;
            9'd170: cos_value = -64540;
            9'd171: cos_value = -64729;
            9'd172: cos_value = -64898;
            9'd173: cos_value = -65047;
            9'd174: cos_value = -65176;
            9'd175: cos_value = -65286;
            9'd176: cos_value = -65376;
            9'd177: cos_value = -65446;
            9'd178: cos_value = -65496;
            9'd179: cos_value = -65526;
            9'd180: cos_value = -65536;
            9'd181: cos_value = -65526;
            9'd182: cos_value = -65496;
            9'd183: cos_value = -65446;
            9'd184: cos_value = -65376;
            9'd185: cos_value = -65286;
            9'd186: cos_value = -65176;
            9'd187: cos_value = -65047;
            9'd188: cos_value = -64898;
            9'd189: cos_value = -64729;
            9'd190: cos_value = -64540;
            9'd191: cos_value = -64331;
            9'd192: cos_value = -64103;
            9'd193: cos_value = -63856;
            9'd194: cos_value = -63589;
            9'd195: cos_value = -63302;
            9'd196: cos_value = -62997;
            9'd197: cos_value = -62672;
            9'd198: cos_value = -62328;
            9'd199: cos_value = -61965;
            9'd200: cos_value = -61583;
            9'd201: cos_value = -61183;
            9'd202: cos_value = -60763;
            9'd203: cos_value = -60326;
            9'd204: cos_value = -59870;
            9'd205: cos_value = -59395;
            9'd206: cos_value = -58903;
            9'd207: cos_value = -58393;
            9'd208: cos_value = -57864;
            9'd209: cos_value = -57319;
            9'd210: cos_value = -56755;
            9'd211: cos_value = -56175;
            9'd212: cos_value = -55577;
            9'd213: cos_value = -54963;
            9'd214: cos_value = -54331;
            9'd215: cos_value = -53683;
            9'd216: cos_value = -53019;
            9'd217: cos_value = -52339;
            9'd218: cos_value = -51643;
            9'd219: cos_value = -50931;
            9'd220: cos_value = -50203;
            9'd221: cos_value = -49460;
            9'd222: cos_value = -48702;
            9'd223: cos_value = -47929;
            9'd224: cos_value = -47142;
            9'd225: cos_value = -46340;
            9'd226: cos_value = -45525;
            9'd227: cos_value = -44695;
            9'd228: cos_value = -43852;
            9'd229: cos_value = -42995;
            9'd230: cos_value = -42125;
            9'd231: cos_value = -41243;
            9'd232: cos_value = -40347;
            9'd233: cos_value = -39440;
            9'd234: cos_value = -38521;
            9'd235: cos_value = -37589;
            9'd236: cos_value = -36647;
            9'd237: cos_value = -35693;
            9'd238: cos_value = -34728;
            9'd239: cos_value = -33753;
            9'd240: cos_value = -32768;
            9'd241: cos_value = -31772;
            9'd242: cos_value = -30767;
            9'd243: cos_value = -29752;
            9'd244: cos_value = -28729;
            9'd245: cos_value = -27696;
            9'd246: cos_value = -26655;
            9'd247: cos_value = -25606;
            9'd248: cos_value = -24550;
            9'd249: cos_value = -23486;
            9'd250: cos_value = -22414;
            9'd251: cos_value = -21336;
            9'd252: cos_value = -20251;
            9'd253: cos_value = -19160;
            9'd254: cos_value = -18064;
            9'd255: cos_value = -16961;
            9'd256: cos_value = -15854;
            9'd257: cos_value = -14742;
            9'd258: cos_value = -13625;
            9'd259: cos_value = -12504;
            9'd260: cos_value = -11380;
            9'd261: cos_value = -10252;
            9'd262: cos_value = -9120;
            9'd263: cos_value = -7986;
            9'd264: cos_value = -6850;
            9'd265: cos_value = -5711;
            9'd266: cos_value = -4571;
            9'd267: cos_value = -3429;
            9'd268: cos_value = -2287;
            9'd269: cos_value = -1143;
            9'd270: cos_value = 0;
            9'd271: cos_value = 1143;
            9'd272: cos_value = 2287;
            9'd273: cos_value = 3429;
            9'd274: cos_value = 4571;
            9'd275: cos_value = 5711;
            9'd276: cos_value = 6850;
            9'd277: cos_value = 7986;
            9'd278: cos_value = 9120;
            9'd279: cos_value = 10252;
            9'd280: cos_value = 11380;
            9'd281: cos_value = 12504;
            9'd282: cos_value = 13625;
            9'd283: cos_value = 14742;
            9'd284: cos_value = 15854;
            9'd285: cos_value = 16961;
            9'd286: cos_value = 18064;
            9'd287: cos_value = 19160;
            9'd288: cos_value = 20251;
            9'd289: cos_value = 21336;
            9'd290: cos_value = 22414;
            9'd291: cos_value = 23486;
            9'd292: cos_value = 24550;
            9'd293: cos_value = 25606;
            9'd294: cos_value = 26655;
            9'd295: cos_value = 27696;
            9'd296: cos_value = 28729;
            9'd297: cos_value = 29752;
            9'd298: cos_value = 30767;
            9'd299: cos_value = 31772;
            9'd300: cos_value = 32768;
            9'd301: cos_value = 33753;
            9'd302: cos_value = 34728;
            9'd303: cos_value = 35693;
            9'd304: cos_value = 36647;
            9'd305: cos_value = 37589;
            9'd306: cos_value = 38521;
            9'd307: cos_value = 39440;
            9'd308: cos_value = 40347;
            9'd309: cos_value = 41243;
            9'd310: cos_value = 42125;
            9'd311: cos_value = 42995;
            9'd312: cos_value = 43852;
            9'd313: cos_value = 44695;
            9'd314: cos_value = 45525;
            9'd315: cos_value = 46340;
            9'd316: cos_value = 47142;
            9'd317: cos_value = 47929;
            9'd318: cos_value = 48702;
            9'd319: cos_value = 49460;
            9'd320: cos_value = 50203;
            9'd321: cos_value = 50931;
            9'd322: cos_value = 51643;
            9'd323: cos_value = 52339;
            9'd324: cos_value = 53019;
            9'd325: cos_value = 53683;
            9'd326: cos_value = 54331;
            9'd327: cos_value = 54963;
            9'd328: cos_value = 55577;
            9'd329: cos_value = 56175;
            9'd330: cos_value = 56755;
            9'd331: cos_value = 57319;
            9'd332: cos_value = 57864;
            9'd333: cos_value = 58393;
            9'd334: cos_value = 58903;
            9'd335: cos_value = 59395;
            9'd336: cos_value = 59870;
            9'd337: cos_value = 60326;
            9'd338: cos_value = 60763;
            9'd339: cos_value = 61183;
            9'd340: cos_value = 61583;
            9'd341: cos_value = 61965;
            9'd342: cos_value = 62328;
            9'd343: cos_value = 62672;
            9'd344: cos_value = 62997;
            9'd345: cos_value = 63302;
            9'd346: cos_value = 63589;
            9'd347: cos_value = 63856;
            9'd348: cos_value = 64103;
            9'd349: cos_value = 64331;
            9'd350: cos_value = 64540;
            9'd351: cos_value = 64729;
            9'd352: cos_value = 64898;
            9'd353: cos_value = 65047;
            9'd354: cos_value = 65176;
            9'd355: cos_value = 65286;
            9'd356: cos_value = 65376;
            9'd357: cos_value = 65446;
            9'd358: cos_value = 65496;
            9'd359: cos_value = 65526;
            default: cos_value = 0;
        endcase
    end
endmodule
