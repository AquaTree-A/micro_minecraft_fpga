module p_transformation (
	input logic x,
	input logic y,
	input logic z,

	output logic x_,
	output logic y_
);
	
	

endmodule