module texture_rom(
    input  logic clk,
    input  logic [4:0] id,
    input  logic [3:0] x,
    input  logic [3:0] y,
    output logic [7:0] data
);

    parameter ADDR_WIDTH = 8;
    parameter DATA_WIDTH = 8;
    parameter TYPE_NUMBER = 22;
    // ROM definition
    parameter [0:22*2**ADDR_WIDTH-1][DATA_WIDTH-1:0] TEXTURE_ROM = {
        // 00_dirt
        8'b00000010, // Color (11, 8, 5) (0, 0)
        8'b00000100, // Color (9, 6, 4) (1, 0)
        8'b00000100, // Color (9, 6, 4) (2, 0)
        8'b00000110, // Color (7, 5, 3) (3, 0)
        8'b00000110, // Color (7, 5, 3) (4, 0)
        8'b00000010, // Color (11, 8, 5) (5, 0)
        8'b00000100, // Color (9, 6, 4) (6, 0)
        8'b00000100, // Color (9, 6, 4) (7, 0)
        8'b00000110, // Color (7, 5, 3) (8, 0)
        8'b00000110, // Color (7, 5, 3) (9, 0)
        8'b00001000, // Color (5, 3, 2) (10, 0)
        8'b00000110, // Color (7, 5, 3) (11, 0)
        8'b00000110, // Color (7, 5, 3) (12, 0)
        8'b00000010, // Color (11, 8, 5) (13, 0)
        8'b00000110, // Color (7, 5, 3) (14, 0)
        8'b00000010, // Color (11, 8, 5) (15, 0)
        8'b00000110, // Color (7, 5, 3) (0, 1)
        8'b00000100, // Color (9, 6, 4) (1, 1)
        8'b00001000, // Color (5, 3, 2) (2, 1)
        8'b00000110, // Color (7, 5, 3) (3, 1)
        8'b00000110, // Color (7, 5, 3) (4, 1)
        8'b00000100, // Color (9, 6, 4) (5, 1)
        8'b00001010, // Color (8, 8, 8) (6, 1)
        8'b00001000, // Color (5, 3, 2) (7, 1)
        8'b00000110, // Color (7, 5, 3) (8, 1)
        8'b00000010, // Color (11, 8, 5) (9, 1)
        8'b00000100, // Color (9, 6, 4) (10, 1)
        8'b00000110, // Color (7, 5, 3) (11, 1)
        8'b00000010, // Color (11, 8, 5) (12, 1)
        8'b00000100, // Color (9, 6, 4) (13, 1)
        8'b00001000, // Color (5, 3, 2) (14, 1)
        8'b00001000, // Color (5, 3, 2) (15, 1)
        8'b00000010, // Color (11, 8, 5) (0, 2)
        8'b00000110, // Color (7, 5, 3) (1, 2)
        8'b00000110, // Color (7, 5, 3) (2, 2)
        8'b00001000, // Color (5, 3, 2) (3, 2)
        8'b00000010, // Color (11, 8, 5) (4, 2)
        8'b00000110, // Color (7, 5, 3) (5, 2)
        8'b00000110, // Color (7, 5, 3) (6, 2)
        8'b00000110, // Color (7, 5, 3) (7, 2)
        8'b00000010, // Color (11, 8, 5) (8, 2)
        8'b00000110, // Color (7, 5, 3) (9, 2)
        8'b00000110, // Color (7, 5, 3) (10, 2)
        8'b00000110, // Color (7, 5, 3) (11, 2)
        8'b00001000, // Color (5, 3, 2) (12, 2)
        8'b00001000, // Color (5, 3, 2) (13, 2)
        8'b00000010, // Color (11, 8, 5) (14, 2)
        8'b00000110, // Color (7, 5, 3) (15, 2)
        8'b00000100, // Color (9, 6, 4) (0, 3)
        8'b00001100, // Color (6, 6, 6) (1, 3)
        8'b00000010, // Color (11, 8, 5) (2, 3)
        8'b00000110, // Color (7, 5, 3) (3, 3)
        8'b00000100, // Color (9, 6, 4) (4, 3)
        8'b00001000, // Color (5, 3, 2) (5, 3)
        8'b00000110, // Color (7, 5, 3) (6, 3)
        8'b00000010, // Color (11, 8, 5) (7, 3)
        8'b00000100, // Color (9, 6, 4) (8, 3)
        8'b00000100, // Color (9, 6, 4) (9, 3)
        8'b00000110, // Color (7, 5, 3) (10, 3)
        8'b00000100, // Color (9, 6, 4) (11, 3)
        8'b00000110, // Color (7, 5, 3) (12, 3)
        8'b00000010, // Color (11, 8, 5) (13, 3)
        8'b00000100, // Color (9, 6, 4) (14, 3)
        8'b00000110, // Color (7, 5, 3) (15, 3)
        8'b00000100, // Color (9, 6, 4) (0, 4)
        8'b00000110, // Color (7, 5, 3) (1, 4)
        8'b00000100, // Color (9, 6, 4) (2, 4)
        8'b00000010, // Color (11, 8, 5) (3, 4)
        8'b00001000, // Color (5, 3, 2) (4, 4)
        8'b00000100, // Color (9, 6, 4) (5, 4)
        8'b00000110, // Color (7, 5, 3) (6, 4)
        8'b00000110, // Color (7, 5, 3) (7, 4)
        8'b00000100, // Color (9, 6, 4) (8, 4)
        8'b00001000, // Color (5, 3, 2) (9, 4)
        8'b00000110, // Color (7, 5, 3) (10, 4)
        8'b00001100, // Color (6, 6, 6) (11, 4)
        8'b00000110, // Color (7, 5, 3) (12, 4)
        8'b00000100, // Color (9, 6, 4) (13, 4)
        8'b00001000, // Color (5, 3, 2) (14, 4)
        8'b00000110, // Color (7, 5, 3) (15, 4)
        8'b00000110, // Color (7, 5, 3) (0, 5)
        8'b00001000, // Color (5, 3, 2) (1, 5)
        8'b00000100, // Color (9, 6, 4) (2, 5)
        8'b00000100, // Color (9, 6, 4) (3, 5)
        8'b00000110, // Color (7, 5, 3) (4, 5)
        8'b00000100, // Color (9, 6, 4) (5, 5)
        8'b00001000, // Color (5, 3, 2) (6, 5)
        8'b00001000, // Color (5, 3, 2) (7, 5)
        8'b00001000, // Color (5, 3, 2) (8, 5)
        8'b00000110, // Color (7, 5, 3) (9, 5)
        8'b00000110, // Color (7, 5, 3) (10, 5)
        8'b00001000, // Color (5, 3, 2) (11, 5)
        8'b00000110, // Color (7, 5, 3) (12, 5)
        8'b00000110, // Color (7, 5, 3) (13, 5)
        8'b00000110, // Color (7, 5, 3) (14, 5)
        8'b00000010, // Color (11, 8, 5) (15, 5)
        8'b00000010, // Color (11, 8, 5) (0, 6)
        8'b00000110, // Color (7, 5, 3) (1, 6)
        8'b00000110, // Color (7, 5, 3) (2, 6)
        8'b00000110, // Color (7, 5, 3) (3, 6)
        8'b00001010, // Color (8, 8, 8) (4, 6)
        8'b00000110, // Color (7, 5, 3) (5, 6)
        8'b00000110, // Color (7, 5, 3) (6, 6)
        8'b00000010, // Color (11, 8, 5) (7, 6)
        8'b00000010, // Color (11, 8, 5) (8, 6)
        8'b00000110, // Color (7, 5, 3) (9, 6)
        8'b00000010, // Color (11, 8, 5) (10, 6)
        8'b00000010, // Color (11, 8, 5) (11, 6)
        8'b00000110, // Color (7, 5, 3) (12, 6)
        8'b00000100, // Color (9, 6, 4) (13, 6)
        8'b00000110, // Color (7, 5, 3) (14, 6)
        8'b00000100, // Color (9, 6, 4) (15, 6)
        8'b00000110, // Color (7, 5, 3) (0, 7)
        8'b00000110, // Color (7, 5, 3) (1, 7)
        8'b00000010, // Color (11, 8, 5) (2, 7)
        8'b00000010, // Color (11, 8, 5) (3, 7)
        8'b00000100, // Color (9, 6, 4) (4, 7)
        8'b00000100, // Color (9, 6, 4) (5, 7)
        8'b00000110, // Color (7, 5, 3) (6, 7)
        8'b00000110, // Color (7, 5, 3) (7, 7)
        8'b00000100, // Color (9, 6, 4) (8, 7)
        8'b00001000, // Color (5, 3, 2) (9, 7)
        8'b00000100, // Color (9, 6, 4) (10, 7)
        8'b00000100, // Color (9, 6, 4) (11, 7)
        8'b00000110, // Color (7, 5, 3) (12, 7)
        8'b00000110, // Color (7, 5, 3) (13, 7)
        8'b00000100, // Color (9, 6, 4) (14, 7)
        8'b00000100, // Color (9, 6, 4) (15, 7)
        8'b00000100, // Color (9, 6, 4) (0, 8)
        8'b00000110, // Color (7, 5, 3) (1, 8)
        8'b00000110, // Color (7, 5, 3) (2, 8)
        8'b00000100, // Color (9, 6, 4) (3, 8)
        8'b00000110, // Color (7, 5, 3) (4, 8)
        8'b00000100, // Color (9, 6, 4) (5, 8)
        8'b00000110, // Color (7, 5, 3) (6, 8)
        8'b00001000, // Color (5, 3, 2) (7, 8)
        8'b00000110, // Color (7, 5, 3) (8, 8)
        8'b00000100, // Color (9, 6, 4) (9, 8)
        8'b00000100, // Color (9, 6, 4) (10, 8)
        8'b00000110, // Color (7, 5, 3) (11, 8)
        8'b00000110, // Color (7, 5, 3) (12, 8)
        8'b00000110, // Color (7, 5, 3) (13, 8)
        8'b00001000, // Color (5, 3, 2) (14, 8)
        8'b00000110, // Color (7, 5, 3) (15, 8)
        8'b00000110, // Color (7, 5, 3) (0, 9)
        8'b00000100, // Color (9, 6, 4) (1, 9)
        8'b00001000, // Color (5, 3, 2) (2, 9)
        8'b00000110, // Color (7, 5, 3) (3, 9)
        8'b00000110, // Color (7, 5, 3) (4, 9)
        8'b00001000, // Color (5, 3, 2) (5, 9)
        8'b00001000, // Color (5, 3, 2) (6, 9)
        8'b00000110, // Color (7, 5, 3) (7, 9)
        8'b00000110, // Color (7, 5, 3) (8, 9)
        8'b00000110, // Color (7, 5, 3) (9, 9)
        8'b00000110, // Color (7, 5, 3) (10, 9)
        8'b00000110, // Color (7, 5, 3) (11, 9)
        8'b00000010, // Color (11, 8, 5) (12, 9)
        8'b00000010, // Color (11, 8, 5) (13, 9)
        8'b00000110, // Color (7, 5, 3) (14, 9)
        8'b00000100, // Color (9, 6, 4) (15, 9)
        8'b00000110, // Color (7, 5, 3) (0, 10)
        8'b00000100, // Color (9, 6, 4) (1, 10)
        8'b00000110, // Color (7, 5, 3) (2, 10)
        8'b00000010, // Color (11, 8, 5) (3, 10)
        8'b00000010, // Color (11, 8, 5) (4, 10)
        8'b00000110, // Color (7, 5, 3) (5, 10)
        8'b00000010, // Color (11, 8, 5) (6, 10)
        8'b00000100, // Color (9, 6, 4) (7, 10)
        8'b00001000, // Color (5, 3, 2) (8, 10)
        8'b00000010, // Color (11, 8, 5) (9, 10)
        8'b00000010, // Color (11, 8, 5) (10, 10)
        8'b00001000, // Color (5, 3, 2) (11, 10)
        8'b00000100, // Color (9, 6, 4) (12, 10)
        8'b00000100, // Color (9, 6, 4) (13, 10)
        8'b00001010, // Color (8, 8, 8) (14, 10)
        8'b00000110, // Color (7, 5, 3) (15, 10)
        8'b00000100, // Color (9, 6, 4) (0, 11)
        8'b00000110, // Color (7, 5, 3) (1, 11)
        8'b00000110, // Color (7, 5, 3) (2, 11)
        8'b00000100, // Color (9, 6, 4) (3, 11)
        8'b00000100, // Color (9, 6, 4) (4, 11)
        8'b00000010, // Color (11, 8, 5) (5, 11)
        8'b00000110, // Color (7, 5, 3) (6, 11)
        8'b00000100, // Color (9, 6, 4) (7, 11)
        8'b00001100, // Color (6, 6, 6) (8, 11)
        8'b00000100, // Color (9, 6, 4) (9, 11)
        8'b00000100, // Color (9, 6, 4) (10, 11)
        8'b00000110, // Color (7, 5, 3) (11, 11)
        8'b00001000, // Color (5, 3, 2) (12, 11)
        8'b00000100, // Color (9, 6, 4) (13, 11)
        8'b00000110, // Color (7, 5, 3) (14, 11)
        8'b00001000, // Color (5, 3, 2) (15, 11)
        8'b00000110, // Color (7, 5, 3) (0, 12)
        8'b00001000, // Color (5, 3, 2) (1, 12)
        8'b00000100, // Color (9, 6, 4) (2, 12)
        8'b00000110, // Color (7, 5, 3) (3, 12)
        8'b00000100, // Color (9, 6, 4) (4, 12)
        8'b00000100, // Color (9, 6, 4) (5, 12)
        8'b00000010, // Color (11, 8, 5) (6, 12)
        8'b00000110, // Color (7, 5, 3) (7, 12)
        8'b00000110, // Color (7, 5, 3) (8, 12)
        8'b00000110, // Color (7, 5, 3) (9, 12)
        8'b00000110, // Color (7, 5, 3) (10, 12)
        8'b00000110, // Color (7, 5, 3) (11, 12)
        8'b00000110, // Color (7, 5, 3) (12, 12)
        8'b00000110, // Color (7, 5, 3) (13, 12)
        8'b00000010, // Color (11, 8, 5) (14, 12)
        8'b00000010, // Color (11, 8, 5) (15, 12)
        8'b00000110, // Color (7, 5, 3) (0, 13)
        8'b00000100, // Color (9, 6, 4) (1, 13)
        8'b00000110, // Color (7, 5, 3) (2, 13)
        8'b00000110, // Color (7, 5, 3) (3, 13)
        8'b00001110, // Color (7, 5, 4) (4, 13)
        8'b00000110, // Color (7, 5, 3) (5, 13)
        8'b00000100, // Color (9, 6, 4) (6, 13)
        8'b00000100, // Color (9, 6, 4) (7, 13)
        8'b00000110, // Color (7, 5, 3) (8, 13)
        8'b00001000, // Color (5, 3, 2) (9, 13)
        8'b00000010, // Color (11, 8, 5) (10, 13)
        8'b00001000, // Color (5, 3, 2) (11, 13)
        8'b00000110, // Color (7, 5, 3) (12, 13)
        8'b00000010, // Color (11, 8, 5) (13, 13)
        8'b00000100, // Color (9, 6, 4) (14, 13)
        8'b00000100, // Color (9, 6, 4) (15, 13)
        8'b00000100, // Color (9, 6, 4) (0, 14)
        8'b00000110, // Color (7, 5, 3) (1, 14)
        8'b00001000, // Color (5, 3, 2) (2, 14)
        8'b00000010, // Color (11, 8, 5) (3, 14)
        8'b00000110, // Color (7, 5, 3) (4, 14)
        8'b00001000, // Color (5, 3, 2) (5, 14)
        8'b00000110, // Color (7, 5, 3) (6, 14)
        8'b00001000, // Color (5, 3, 2) (7, 14)
        8'b00000010, // Color (11, 8, 5) (8, 14)
        8'b00000010, // Color (11, 8, 5) (9, 14)
        8'b00000110, // Color (7, 5, 3) (10, 14)
        8'b00000100, // Color (9, 6, 4) (11, 14)
        8'b00000110, // Color (7, 5, 3) (12, 14)
        8'b00000110, // Color (7, 5, 3) (13, 14)
        8'b00000100, // Color (9, 6, 4) (14, 14)
        8'b00000100, // Color (9, 6, 4) (15, 14)
        8'b00000100, // Color (9, 6, 4) (0, 15)
        8'b00000110, // Color (7, 5, 3) (1, 15)
        8'b00000010, // Color (11, 8, 5) (2, 15)
        8'b00000100, // Color (9, 6, 4) (3, 15)
        8'b00000100, // Color (9, 6, 4) (4, 15)
        8'b00000110, // Color (7, 5, 3) (5, 15)
        8'b00001010, // Color (8, 8, 8) (6, 15)
        8'b00000110, // Color (7, 5, 3) (7, 15)
        8'b00000100, // Color (9, 6, 4) (8, 15)
        8'b00000100, // Color (9, 6, 4) (9, 15)
        8'b00000110, // Color (7, 5, 3) (10, 15)
        8'b00000110, // Color (7, 5, 3) (11, 15)
        8'b00000100, // Color (9, 6, 4) (12, 15)
        8'b00000100, // Color (9, 6, 4) (13, 15)
        8'b00000110, // Color (7, 5, 3) (14, 15)
        8'b00001000, // Color (5, 3, 2) (15, 15)
        // 01_grass_side
        8'b00010000, // Color (7, 11, 4) (0, 0)
        8'b00010000, // Color (7, 11, 4) (1, 0)
        8'b00010000, // Color (7, 11, 4) (2, 0)
        8'b00010010, // Color (6, 10, 3) (3, 0)
        8'b00010010, // Color (6, 10, 3) (4, 0)
        8'b00010100, // Color (6, 10, 4) (5, 0)
        8'b00010110, // Color (5, 9, 3) (6, 0)
        8'b00010100, // Color (6, 10, 4) (7, 0)
        8'b00011000, // Color (7, 11, 5) (8, 0)
        8'b00010000, // Color (7, 11, 4) (9, 0)
        8'b00010100, // Color (6, 10, 4) (10, 0)
        8'b00010010, // Color (6, 10, 3) (11, 0)
        8'b00010010, // Color (6, 10, 3) (12, 0)
        8'b00010010, // Color (6, 10, 3) (13, 0)
        8'b00011010, // Color (5, 9, 2) (14, 0)
        8'b00010100, // Color (6, 10, 4) (15, 0)
        8'b00010000, // Color (7, 11, 4) (0, 1)
        8'b00010100, // Color (6, 10, 4) (1, 1)
        8'b00011100, // Color (8, 11, 5) (2, 1)
        8'b00011100, // Color (8, 11, 5) (3, 1)
        8'b00011100, // Color (8, 11, 5) (4, 1)
        8'b00001000, // Color (5, 3, 2) (5, 1)
        8'b00010010, // Color (6, 10, 3) (6, 1)
        8'b00010010, // Color (6, 10, 3) (7, 1)
        8'b00010110, // Color (5, 9, 3) (8, 1)
        8'b00011110, // Color (9, 12, 6) (9, 1)
        8'b00100000, // Color (9, 11, 6) (10, 1)
        8'b00010000, // Color (7, 11, 4) (11, 1)
        8'b00010010, // Color (6, 10, 3) (12, 1)
        8'b00010100, // Color (6, 10, 4) (13, 1)
        8'b00010010, // Color (6, 10, 3) (14, 1)
        8'b00010100, // Color (6, 10, 4) (15, 1)
        8'b00011100, // Color (8, 11, 5) (0, 2)
        8'b00001000, // Color (5, 3, 2) (1, 2)
        8'b00011110, // Color (9, 12, 6) (2, 2)
        8'b00010010, // Color (6, 10, 3) (3, 2)
        8'b00010010, // Color (6, 10, 3) (4, 2)
        8'b00001000, // Color (5, 3, 2) (5, 2)
        8'b00010000, // Color (7, 11, 4) (6, 2)
        8'b00001000, // Color (5, 3, 2) (7, 2)
        8'b00010000, // Color (7, 11, 4) (8, 2)
        8'b00011000, // Color (7, 11, 5) (9, 2)
        8'b00011110, // Color (9, 12, 6) (10, 2)
        8'b00011110, // Color (9, 12, 6) (11, 2)
        8'b00001000, // Color (5, 3, 2) (12, 2)
        8'b00011010, // Color (5, 9, 2) (13, 2)
        8'b00010010, // Color (6, 10, 3) (14, 2)
        8'b00001000, // Color (5, 3, 2) (15, 2)
        8'b00001000, // Color (5, 3, 2) (0, 3)
        8'b00001100, // Color (6, 6, 6) (1, 3)
        8'b00001000, // Color (5, 3, 2) (2, 3)
        8'b00001000, // Color (5, 3, 2) (3, 3)
        8'b00010000, // Color (7, 11, 4) (4, 3)
        8'b00001000, // Color (5, 3, 2) (5, 3)
        8'b00001000, // Color (5, 3, 2) (6, 3)
        8'b00001000, // Color (5, 3, 2) (7, 3)
        8'b00010110, // Color (5, 9, 3) (8, 3)
        8'b00001000, // Color (5, 3, 2) (9, 3)
        8'b00010100, // Color (6, 10, 4) (10, 3)
        8'b00001000, // Color (5, 3, 2) (11, 3)
        8'b00000110, // Color (7, 5, 3) (12, 3)
        8'b00001000, // Color (5, 3, 2) (13, 3)
        8'b00001000, // Color (5, 3, 2) (14, 3)
        8'b00000110, // Color (7, 5, 3) (15, 3)
        8'b00000100, // Color (9, 6, 4) (0, 4)
        8'b00000110, // Color (7, 5, 3) (1, 4)
        8'b00000100, // Color (9, 6, 4) (2, 4)
        8'b00000010, // Color (11, 8, 5) (3, 4)
        8'b00001000, // Color (5, 3, 2) (4, 4)
        8'b00000100, // Color (9, 6, 4) (5, 4)
        8'b00000110, // Color (7, 5, 3) (6, 4)
        8'b00000110, // Color (7, 5, 3) (7, 4)
        8'b00001000, // Color (5, 3, 2) (8, 4)
        8'b00001000, // Color (5, 3, 2) (9, 4)
        8'b00001000, // Color (5, 3, 2) (10, 4)
        8'b00001100, // Color (6, 6, 6) (11, 4)
        8'b00000110, // Color (7, 5, 3) (12, 4)
        8'b00000100, // Color (9, 6, 4) (13, 4)
        8'b00001000, // Color (5, 3, 2) (14, 4)
        8'b00000110, // Color (7, 5, 3) (15, 4)
        8'b00000110, // Color (7, 5, 3) (0, 5)
        8'b00001000, // Color (5, 3, 2) (1, 5)
        8'b00000100, // Color (9, 6, 4) (2, 5)
        8'b00000100, // Color (9, 6, 4) (3, 5)
        8'b00000110, // Color (7, 5, 3) (4, 5)
        8'b00000100, // Color (9, 6, 4) (5, 5)
        8'b00001000, // Color (5, 3, 2) (6, 5)
        8'b00001000, // Color (5, 3, 2) (7, 5)
        8'b00001000, // Color (5, 3, 2) (8, 5)
        8'b00000110, // Color (7, 5, 3) (9, 5)
        8'b00000110, // Color (7, 5, 3) (10, 5)
        8'b00001000, // Color (5, 3, 2) (11, 5)
        8'b00000110, // Color (7, 5, 3) (12, 5)
        8'b00000110, // Color (7, 5, 3) (13, 5)
        8'b00000110, // Color (7, 5, 3) (14, 5)
        8'b00000010, // Color (11, 8, 5) (15, 5)
        8'b00000010, // Color (11, 8, 5) (0, 6)
        8'b00000110, // Color (7, 5, 3) (1, 6)
        8'b00000110, // Color (7, 5, 3) (2, 6)
        8'b00000110, // Color (7, 5, 3) (3, 6)
        8'b00001010, // Color (8, 8, 8) (4, 6)
        8'b00000110, // Color (7, 5, 3) (5, 6)
        8'b00000110, // Color (7, 5, 3) (6, 6)
        8'b00000010, // Color (11, 8, 5) (7, 6)
        8'b00000010, // Color (11, 8, 5) (8, 6)
        8'b00000110, // Color (7, 5, 3) (9, 6)
        8'b00000010, // Color (11, 8, 5) (10, 6)
        8'b00000010, // Color (11, 8, 5) (11, 6)
        8'b00000110, // Color (7, 5, 3) (12, 6)
        8'b00000100, // Color (9, 6, 4) (13, 6)
        8'b00000110, // Color (7, 5, 3) (14, 6)
        8'b00000100, // Color (9, 6, 4) (15, 6)
        8'b00000110, // Color (7, 5, 3) (0, 7)
        8'b00000110, // Color (7, 5, 3) (1, 7)
        8'b00000010, // Color (11, 8, 5) (2, 7)
        8'b00000010, // Color (11, 8, 5) (3, 7)
        8'b00000100, // Color (9, 6, 4) (4, 7)
        8'b00000100, // Color (9, 6, 4) (5, 7)
        8'b00000110, // Color (7, 5, 3) (6, 7)
        8'b00000110, // Color (7, 5, 3) (7, 7)
        8'b00000100, // Color (9, 6, 4) (8, 7)
        8'b00001000, // Color (5, 3, 2) (9, 7)
        8'b00000100, // Color (9, 6, 4) (10, 7)
        8'b00000100, // Color (9, 6, 4) (11, 7)
        8'b00000110, // Color (7, 5, 3) (12, 7)
        8'b00000110, // Color (7, 5, 3) (13, 7)
        8'b00000100, // Color (9, 6, 4) (14, 7)
        8'b00000100, // Color (9, 6, 4) (15, 7)
        8'b00000100, // Color (9, 6, 4) (0, 8)
        8'b00000110, // Color (7, 5, 3) (1, 8)
        8'b00000110, // Color (7, 5, 3) (2, 8)
        8'b00000100, // Color (9, 6, 4) (3, 8)
        8'b00000110, // Color (7, 5, 3) (4, 8)
        8'b00000100, // Color (9, 6, 4) (5, 8)
        8'b00000110, // Color (7, 5, 3) (6, 8)
        8'b00001000, // Color (5, 3, 2) (7, 8)
        8'b00000110, // Color (7, 5, 3) (8, 8)
        8'b00000100, // Color (9, 6, 4) (9, 8)
        8'b00000100, // Color (9, 6, 4) (10, 8)
        8'b00000110, // Color (7, 5, 3) (11, 8)
        8'b00000110, // Color (7, 5, 3) (12, 8)
        8'b00000110, // Color (7, 5, 3) (13, 8)
        8'b00001000, // Color (5, 3, 2) (14, 8)
        8'b00000110, // Color (7, 5, 3) (15, 8)
        8'b00000110, // Color (7, 5, 3) (0, 9)
        8'b00000100, // Color (9, 6, 4) (1, 9)
        8'b00001000, // Color (5, 3, 2) (2, 9)
        8'b00000110, // Color (7, 5, 3) (3, 9)
        8'b00000110, // Color (7, 5, 3) (4, 9)
        8'b00001000, // Color (5, 3, 2) (5, 9)
        8'b00001000, // Color (5, 3, 2) (6, 9)
        8'b00000110, // Color (7, 5, 3) (7, 9)
        8'b00000110, // Color (7, 5, 3) (8, 9)
        8'b00000110, // Color (7, 5, 3) (9, 9)
        8'b00000110, // Color (7, 5, 3) (10, 9)
        8'b00000110, // Color (7, 5, 3) (11, 9)
        8'b00000010, // Color (11, 8, 5) (12, 9)
        8'b00000010, // Color (11, 8, 5) (13, 9)
        8'b00000110, // Color (7, 5, 3) (14, 9)
        8'b00000100, // Color (9, 6, 4) (15, 9)
        8'b00000110, // Color (7, 5, 3) (0, 10)
        8'b00000100, // Color (9, 6, 4) (1, 10)
        8'b00000110, // Color (7, 5, 3) (2, 10)
        8'b00000010, // Color (11, 8, 5) (3, 10)
        8'b00000010, // Color (11, 8, 5) (4, 10)
        8'b00000110, // Color (7, 5, 3) (5, 10)
        8'b00000010, // Color (11, 8, 5) (6, 10)
        8'b00000100, // Color (9, 6, 4) (7, 10)
        8'b00001000, // Color (5, 3, 2) (8, 10)
        8'b00000010, // Color (11, 8, 5) (9, 10)
        8'b00000010, // Color (11, 8, 5) (10, 10)
        8'b00001000, // Color (5, 3, 2) (11, 10)
        8'b00000100, // Color (9, 6, 4) (12, 10)
        8'b00000100, // Color (9, 6, 4) (13, 10)
        8'b00001010, // Color (8, 8, 8) (14, 10)
        8'b00000110, // Color (7, 5, 3) (15, 10)
        8'b00000100, // Color (9, 6, 4) (0, 11)
        8'b00000110, // Color (7, 5, 3) (1, 11)
        8'b00000110, // Color (7, 5, 3) (2, 11)
        8'b00000100, // Color (9, 6, 4) (3, 11)
        8'b00000100, // Color (9, 6, 4) (4, 11)
        8'b00000010, // Color (11, 8, 5) (5, 11)
        8'b00000110, // Color (7, 5, 3) (6, 11)
        8'b00000100, // Color (9, 6, 4) (7, 11)
        8'b00001100, // Color (6, 6, 6) (8, 11)
        8'b00000100, // Color (9, 6, 4) (9, 11)
        8'b00000100, // Color (9, 6, 4) (10, 11)
        8'b00000110, // Color (7, 5, 3) (11, 11)
        8'b00001000, // Color (5, 3, 2) (12, 11)
        8'b00000100, // Color (9, 6, 4) (13, 11)
        8'b00000110, // Color (7, 5, 3) (14, 11)
        8'b00001000, // Color (5, 3, 2) (15, 11)
        8'b00000110, // Color (7, 5, 3) (0, 12)
        8'b00001000, // Color (5, 3, 2) (1, 12)
        8'b00000100, // Color (9, 6, 4) (2, 12)
        8'b00000110, // Color (7, 5, 3) (3, 12)
        8'b00000100, // Color (9, 6, 4) (4, 12)
        8'b00000100, // Color (9, 6, 4) (5, 12)
        8'b00000010, // Color (11, 8, 5) (6, 12)
        8'b00000110, // Color (7, 5, 3) (7, 12)
        8'b00000110, // Color (7, 5, 3) (8, 12)
        8'b00000110, // Color (7, 5, 3) (9, 12)
        8'b00000110, // Color (7, 5, 3) (10, 12)
        8'b00000110, // Color (7, 5, 3) (11, 12)
        8'b00000110, // Color (7, 5, 3) (12, 12)
        8'b00000110, // Color (7, 5, 3) (13, 12)
        8'b00000010, // Color (11, 8, 5) (14, 12)
        8'b00000010, // Color (11, 8, 5) (15, 12)
        8'b00000110, // Color (7, 5, 3) (0, 13)
        8'b00000100, // Color (9, 6, 4) (1, 13)
        8'b00000110, // Color (7, 5, 3) (2, 13)
        8'b00000110, // Color (7, 5, 3) (3, 13)
        8'b00001110, // Color (7, 5, 4) (4, 13)
        8'b00000110, // Color (7, 5, 3) (5, 13)
        8'b00000100, // Color (9, 6, 4) (6, 13)
        8'b00000100, // Color (9, 6, 4) (7, 13)
        8'b00000110, // Color (7, 5, 3) (8, 13)
        8'b00001000, // Color (5, 3, 2) (9, 13)
        8'b00000010, // Color (11, 8, 5) (10, 13)
        8'b00001000, // Color (5, 3, 2) (11, 13)
        8'b00000110, // Color (7, 5, 3) (12, 13)
        8'b00000010, // Color (11, 8, 5) (13, 13)
        8'b00000100, // Color (9, 6, 4) (14, 13)
        8'b00000100, // Color (9, 6, 4) (15, 13)
        8'b00000100, // Color (9, 6, 4) (0, 14)
        8'b00000110, // Color (7, 5, 3) (1, 14)
        8'b00001000, // Color (5, 3, 2) (2, 14)
        8'b00000010, // Color (11, 8, 5) (3, 14)
        8'b00000110, // Color (7, 5, 3) (4, 14)
        8'b00001000, // Color (5, 3, 2) (5, 14)
        8'b00000110, // Color (7, 5, 3) (6, 14)
        8'b00001000, // Color (5, 3, 2) (7, 14)
        8'b00000010, // Color (11, 8, 5) (8, 14)
        8'b00000010, // Color (11, 8, 5) (9, 14)
        8'b00000110, // Color (7, 5, 3) (10, 14)
        8'b00000100, // Color (9, 6, 4) (11, 14)
        8'b00000110, // Color (7, 5, 3) (12, 14)
        8'b00000110, // Color (7, 5, 3) (13, 14)
        8'b00000100, // Color (9, 6, 4) (14, 14)
        8'b00000100, // Color (9, 6, 4) (15, 14)
        8'b00000100, // Color (9, 6, 4) (0, 15)
        8'b00000110, // Color (7, 5, 3) (1, 15)
        8'b00000010, // Color (11, 8, 5) (2, 15)
        8'b00000100, // Color (9, 6, 4) (3, 15)
        8'b00000100, // Color (9, 6, 4) (4, 15)
        8'b00000110, // Color (7, 5, 3) (5, 15)
        8'b00001010, // Color (8, 8, 8) (6, 15)
        8'b00000110, // Color (7, 5, 3) (7, 15)
        8'b00000100, // Color (9, 6, 4) (8, 15)
        8'b00000100, // Color (9, 6, 4) (9, 15)
        8'b00000110, // Color (7, 5, 3) (10, 15)
        8'b00000110, // Color (7, 5, 3) (11, 15)
        8'b00000100, // Color (9, 6, 4) (12, 15)
        8'b00000100, // Color (9, 6, 4) (13, 15)
        8'b00000110, // Color (7, 5, 3) (14, 15)
        8'b00001000, // Color (5, 3, 2) (15, 15)
        // 02_grass_top
        8'b00100010, // Color (6, 9, 3) (0, 0)
        8'b00100100, // Color (8, 12, 4) (1, 0)
        8'b00100010, // Color (6, 9, 3) (2, 0)
        8'b00100110, // Color (5, 8, 3) (3, 0)
        8'b00100110, // Color (5, 8, 3) (4, 0)
        8'b00010110, // Color (5, 9, 3) (5, 0)
        8'b00100110, // Color (5, 8, 3) (6, 0)
        8'b00100110, // Color (5, 8, 3) (7, 0)
        8'b00010010, // Color (6, 10, 3) (8, 0)
        8'b00100010, // Color (6, 9, 3) (9, 0)
        8'b00100110, // Color (5, 8, 3) (10, 0)
        8'b00100110, // Color (5, 8, 3) (11, 0)
        8'b00100110, // Color (5, 8, 3) (12, 0)
        8'b00010100, // Color (6, 10, 4) (13, 0)
        8'b00101000, // Color (4, 7, 2) (14, 0)
        8'b00010110, // Color (5, 9, 3) (15, 0)
        8'b00100010, // Color (6, 9, 3) (0, 1)
        8'b00100110, // Color (5, 8, 3) (1, 1)
        8'b00010100, // Color (6, 10, 4) (2, 1)
        8'b00100010, // Color (6, 9, 3) (3, 1)
        8'b00100010, // Color (6, 9, 3) (4, 1)
        8'b00100110, // Color (5, 8, 3) (5, 1)
        8'b00100010, // Color (6, 9, 3) (6, 1)
        8'b00100110, // Color (5, 8, 3) (7, 1)
        8'b00100110, // Color (5, 8, 3) (8, 1)
        8'b00010100, // Color (6, 10, 4) (9, 1)
        8'b00010100, // Color (6, 10, 4) (10, 1)
        8'b00100010, // Color (6, 9, 3) (11, 1)
        8'b00100100, // Color (8, 12, 4) (12, 1)
        8'b00100110, // Color (5, 8, 3) (13, 1)
        8'b00100110, // Color (5, 8, 3) (14, 1)
        8'b00100110, // Color (5, 8, 3) (15, 1)
        8'b00010100, // Color (6, 10, 4) (0, 2)
        8'b00010110, // Color (5, 9, 3) (1, 2)
        8'b00101010, // Color (5, 7, 3) (2, 2)
        8'b00100110, // Color (5, 8, 3) (3, 2)
        8'b00100110, // Color (5, 8, 3) (4, 2)
        8'b00100110, // Color (5, 8, 3) (5, 2)
        8'b00100010, // Color (6, 9, 3) (6, 2)
        8'b00100010, // Color (6, 9, 3) (7, 2)
        8'b00100010, // Color (6, 9, 3) (8, 2)
        8'b00010010, // Color (6, 10, 3) (9, 2)
        8'b00010100, // Color (6, 10, 4) (10, 2)
        8'b00010000, // Color (7, 11, 4) (11, 2)
        8'b00100110, // Color (5, 8, 3) (12, 2)
        8'b00101100, // Color (4, 7, 3) (13, 2)
        8'b00100110, // Color (5, 8, 3) (14, 2)
        8'b00010000, // Color (7, 11, 4) (15, 2)
        8'b00101100, // Color (4, 7, 3) (0, 3)
        8'b00100110, // Color (5, 8, 3) (1, 3)
        8'b00100110, // Color (5, 8, 3) (2, 3)
        8'b00100010, // Color (6, 9, 3) (3, 3)
        8'b00100010, // Color (6, 9, 3) (4, 3)
        8'b00100010, // Color (6, 9, 3) (5, 3)
        8'b00101010, // Color (5, 7, 3) (6, 3)
        8'b00100010, // Color (6, 9, 3) (7, 3)
        8'b00100110, // Color (5, 8, 3) (8, 3)
        8'b00100110, // Color (5, 8, 3) (9, 3)
        8'b00010110, // Color (5, 9, 3) (10, 3)
        8'b00100010, // Color (6, 9, 3) (11, 3)
        8'b00010110, // Color (5, 9, 3) (12, 3)
        8'b00100110, // Color (5, 8, 3) (13, 3)
        8'b00010100, // Color (6, 10, 4) (14, 3)
        8'b00101010, // Color (5, 7, 3) (15, 3)
        8'b00010100, // Color (6, 10, 4) (0, 4)
        8'b00100110, // Color (5, 8, 3) (1, 4)
        8'b00010000, // Color (7, 11, 4) (2, 4)
        8'b00100110, // Color (5, 8, 3) (3, 4)
        8'b00101110, // Color (7, 10, 4) (4, 4)
        8'b00010000, // Color (7, 11, 4) (5, 4)
        8'b00100110, // Color (5, 8, 3) (6, 4)
        8'b00101110, // Color (7, 10, 4) (7, 4)
        8'b00010000, // Color (7, 11, 4) (8, 4)
        8'b00101000, // Color (4, 7, 2) (9, 4)
        8'b00100110, // Color (5, 8, 3) (10, 4)
        8'b00010100, // Color (6, 10, 4) (11, 4)
        8'b00101110, // Color (7, 10, 4) (12, 4)
        8'b00100110, // Color (5, 8, 3) (13, 4)
        8'b00100110, // Color (5, 8, 3) (14, 4)
        8'b00010110, // Color (5, 9, 3) (15, 4)
        8'b00100010, // Color (6, 9, 3) (0, 5)
        8'b00100010, // Color (6, 9, 3) (1, 5)
        8'b00101100, // Color (4, 7, 3) (2, 5)
        8'b00010100, // Color (6, 10, 4) (3, 5)
        8'b00100110, // Color (5, 8, 3) (4, 5)
        8'b00100010, // Color (6, 9, 3) (5, 5)
        8'b00100010, // Color (6, 9, 3) (6, 5)
        8'b00100010, // Color (6, 9, 3) (7, 5)
        8'b00100110, // Color (5, 8, 3) (8, 5)
        8'b00100010, // Color (6, 9, 3) (9, 5)
        8'b00100110, // Color (5, 8, 3) (10, 5)
        8'b00100110, // Color (5, 8, 3) (11, 5)
        8'b00101100, // Color (4, 7, 3) (12, 5)
        8'b00100110, // Color (5, 8, 3) (13, 5)
        8'b00010110, // Color (5, 9, 3) (14, 5)
        8'b00100010, // Color (6, 9, 3) (15, 5)
        8'b00100110, // Color (5, 8, 3) (0, 6)
        8'b00100010, // Color (6, 9, 3) (1, 6)
        8'b00010100, // Color (6, 10, 4) (2, 6)
        8'b00100010, // Color (6, 9, 3) (3, 6)
        8'b00100010, // Color (6, 9, 3) (4, 6)
        8'b00100110, // Color (5, 8, 3) (5, 6)
        8'b00100110, // Color (5, 8, 3) (6, 6)
        8'b00100110, // Color (5, 8, 3) (7, 6)
        8'b00100110, // Color (5, 8, 3) (8, 6)
        8'b00100110, // Color (5, 8, 3) (9, 6)
        8'b00010000, // Color (7, 11, 4) (10, 6)
        8'b00101110, // Color (7, 10, 4) (11, 6)
        8'b00100010, // Color (6, 9, 3) (12, 6)
        8'b00010100, // Color (6, 10, 4) (13, 6)
        8'b00100010, // Color (6, 9, 3) (14, 6)
        8'b00010110, // Color (5, 9, 3) (15, 6)
        8'b00010110, // Color (5, 9, 3) (0, 7)
        8'b00100110, // Color (5, 8, 3) (1, 7)
        8'b00010010, // Color (6, 10, 3) (2, 7)
        8'b00100110, // Color (5, 8, 3) (3, 7)
        8'b00100010, // Color (6, 9, 3) (4, 7)
        8'b00101010, // Color (5, 7, 3) (5, 7)
        8'b00010100, // Color (6, 10, 4) (6, 7)
        8'b00100110, // Color (5, 8, 3) (7, 7)
        8'b00100010, // Color (6, 9, 3) (8, 7)
        8'b00010000, // Color (7, 11, 4) (9, 7)
        8'b00100110, // Color (5, 8, 3) (10, 7)
        8'b00100110, // Color (5, 8, 3) (11, 7)
        8'b00010110, // Color (5, 9, 3) (12, 7)
        8'b00010100, // Color (6, 10, 4) (13, 7)
        8'b00100110, // Color (5, 8, 3) (14, 7)
        8'b00010100, // Color (6, 10, 4) (15, 7)
        8'b00010100, // Color (6, 10, 4) (0, 8)
        8'b00100010, // Color (6, 9, 3) (1, 8)
        8'b00010000, // Color (7, 11, 4) (2, 8)
        8'b00101110, // Color (7, 10, 4) (3, 8)
        8'b00101110, // Color (7, 10, 4) (4, 8)
        8'b00100110, // Color (5, 8, 3) (5, 8)
        8'b00010000, // Color (7, 11, 4) (6, 8)
        8'b00100010, // Color (6, 9, 3) (7, 8)
        8'b00010000, // Color (7, 11, 4) (8, 8)
        8'b00101110, // Color (7, 10, 4) (9, 8)
        8'b00100110, // Color (5, 8, 3) (10, 8)
        8'b00100010, // Color (6, 9, 3) (11, 8)
        8'b00100110, // Color (5, 8, 3) (12, 8)
        8'b00100010, // Color (6, 9, 3) (13, 8)
        8'b00010010, // Color (6, 10, 3) (14, 8)
        8'b00100110, // Color (5, 8, 3) (15, 8)
        8'b00100010, // Color (6, 9, 3) (0, 9)
        8'b00100110, // Color (5, 8, 3) (1, 9)
        8'b00010000, // Color (7, 11, 4) (2, 9)
        8'b00010110, // Color (5, 9, 3) (3, 9)
        8'b00100110, // Color (5, 8, 3) (4, 9)
        8'b00100010, // Color (6, 9, 3) (5, 9)
        8'b00101110, // Color (7, 10, 4) (6, 9)
        8'b00100110, // Color (5, 8, 3) (7, 9)
        8'b00100110, // Color (5, 8, 3) (8, 9)
        8'b00100010, // Color (6, 9, 3) (9, 9)
        8'b00100010, // Color (6, 9, 3) (10, 9)
        8'b00010100, // Color (6, 10, 4) (11, 9)
        8'b00010110, // Color (5, 9, 3) (12, 9)
        8'b00010000, // Color (7, 11, 4) (13, 9)
        8'b00010110, // Color (5, 9, 3) (14, 9)
        8'b00100110, // Color (5, 8, 3) (15, 9)
        8'b00100010, // Color (6, 9, 3) (0, 10)
        8'b00010010, // Color (6, 10, 3) (1, 10)
        8'b00100010, // Color (6, 9, 3) (2, 10)
        8'b00010100, // Color (6, 10, 4) (3, 10)
        8'b00100110, // Color (5, 8, 3) (4, 10)
        8'b00010000, // Color (7, 11, 4) (5, 10)
        8'b00010110, // Color (5, 9, 3) (6, 10)
        8'b00100010, // Color (6, 9, 3) (7, 10)
        8'b00110000, // Color (7, 12, 4) (8, 10)
        8'b00101010, // Color (5, 7, 3) (9, 10)
        8'b00010100, // Color (6, 10, 4) (10, 10)
        8'b00100110, // Color (5, 8, 3) (11, 10)
        8'b00010110, // Color (5, 9, 3) (12, 10)
        8'b00100110, // Color (5, 8, 3) (13, 10)
        8'b00100010, // Color (6, 9, 3) (14, 10)
        8'b00010110, // Color (5, 9, 3) (15, 10)
        8'b00100110, // Color (5, 8, 3) (0, 11)
        8'b00010000, // Color (7, 11, 4) (1, 11)
        8'b00100110, // Color (5, 8, 3) (2, 11)
        8'b00010100, // Color (6, 10, 4) (3, 11)
        8'b00100010, // Color (6, 9, 3) (4, 11)
        8'b00100110, // Color (5, 8, 3) (5, 11)
        8'b00100010, // Color (6, 9, 3) (6, 11)
        8'b00100110, // Color (5, 8, 3) (7, 11)
        8'b00100010, // Color (6, 9, 3) (8, 11)
        8'b00100010, // Color (6, 9, 3) (9, 11)
        8'b00100110, // Color (5, 8, 3) (10, 11)
        8'b00101010, // Color (5, 7, 3) (11, 11)
        8'b00010000, // Color (7, 11, 4) (12, 11)
        8'b00100110, // Color (5, 8, 3) (13, 11)
        8'b00101010, // Color (5, 7, 3) (14, 11)
        8'b00100110, // Color (5, 8, 3) (15, 11)
        8'b00010000, // Color (7, 11, 4) (0, 12)
        8'b00100010, // Color (6, 9, 3) (1, 12)
        8'b00100110, // Color (5, 8, 3) (2, 12)
        8'b00100110, // Color (5, 8, 3) (3, 12)
        8'b00100010, // Color (6, 9, 3) (4, 12)
        8'b00100010, // Color (6, 9, 3) (5, 12)
        8'b00100110, // Color (5, 8, 3) (6, 12)
        8'b00101010, // Color (5, 7, 3) (7, 12)
        8'b00100110, // Color (5, 8, 3) (8, 12)
        8'b00100010, // Color (6, 9, 3) (9, 12)
        8'b00100110, // Color (5, 8, 3) (10, 12)
        8'b00101010, // Color (5, 7, 3) (11, 12)
        8'b00010010, // Color (6, 10, 3) (12, 12)
        8'b00010100, // Color (6, 10, 4) (13, 12)
        8'b00101010, // Color (5, 7, 3) (14, 12)
        8'b00100010, // Color (6, 9, 3) (15, 12)
        8'b00100110, // Color (5, 8, 3) (0, 13)
        8'b00010100, // Color (6, 10, 4) (1, 13)
        8'b00101100, // Color (4, 7, 3) (2, 13)
        8'b00100010, // Color (6, 9, 3) (3, 13)
        8'b00101010, // Color (5, 7, 3) (4, 13)
        8'b00100010, // Color (6, 9, 3) (5, 13)
        8'b00100110, // Color (5, 8, 3) (6, 13)
        8'b00100100, // Color (8, 12, 4) (7, 13)
        8'b00010100, // Color (6, 10, 4) (8, 13)
        8'b00100010, // Color (6, 9, 3) (9, 13)
        8'b00010100, // Color (6, 10, 4) (10, 13)
        8'b00100010, // Color (6, 9, 3) (11, 13)
        8'b00010100, // Color (6, 10, 4) (12, 13)
        8'b00100110, // Color (5, 8, 3) (13, 13)
        8'b00010100, // Color (6, 10, 4) (14, 13)
        8'b00010000, // Color (7, 11, 4) (15, 13)
        8'b00010100, // Color (6, 10, 4) (0, 14)
        8'b00010100, // Color (6, 10, 4) (1, 14)
        8'b00110000, // Color (7, 12, 4) (2, 14)
        8'b00101010, // Color (5, 7, 3) (3, 14)
        8'b00010000, // Color (7, 11, 4) (4, 14)
        8'b00101110, // Color (7, 10, 4) (5, 14)
        8'b00100010, // Color (6, 9, 3) (6, 14)
        8'b00100010, // Color (6, 9, 3) (7, 14)
        8'b00100110, // Color (5, 8, 3) (8, 14)
        8'b00100010, // Color (6, 9, 3) (9, 14)
        8'b00100010, // Color (6, 9, 3) (10, 14)
        8'b00100110, // Color (5, 8, 3) (11, 14)
        8'b00010100, // Color (6, 10, 4) (12, 14)
        8'b00010010, // Color (6, 10, 3) (13, 14)
        8'b00100110, // Color (5, 8, 3) (14, 14)
        8'b00101010, // Color (5, 7, 3) (15, 14)
        8'b00100110, // Color (5, 8, 3) (0, 15)
        8'b00100010, // Color (6, 9, 3) (1, 15)
        8'b00100110, // Color (5, 8, 3) (2, 15)
        8'b00100110, // Color (5, 8, 3) (3, 15)
        8'b00010100, // Color (6, 10, 4) (4, 15)
        8'b00100010, // Color (6, 9, 3) (5, 15)
        8'b00100010, // Color (6, 9, 3) (6, 15)
        8'b00100010, // Color (6, 9, 3) (7, 15)
        8'b00010110, // Color (5, 9, 3) (8, 15)
        8'b00110000, // Color (7, 12, 4) (9, 15)
        8'b00101010, // Color (5, 7, 3) (10, 15)
        8'b00010100, // Color (6, 10, 4) (11, 15)
        8'b00100110, // Color (5, 8, 3) (12, 15)
        8'b00100010, // Color (6, 9, 3) (13, 15)
        8'b00100110, // Color (5, 8, 3) (14, 15)
        8'b00010010, // Color (6, 10, 3) (15, 15)
        // 03_oak_log
        8'b00000110, // Color (7, 5, 3) (0, 0)
        8'b00110010, // Color (4, 3, 2) (1, 0)
        8'b00110100, // Color (9, 7, 4) (2, 0)
        8'b00000110, // Color (7, 5, 3) (3, 0)
        8'b00000110, // Color (7, 5, 3) (4, 0)
        8'b00110110, // Color (3, 2, 1) (5, 0)
        8'b00110100, // Color (9, 7, 4) (6, 0)
        8'b00000110, // Color (7, 5, 3) (7, 0)
        8'b00000110, // Color (7, 5, 3) (8, 0)
        8'b00110110, // Color (3, 2, 1) (9, 0)
        8'b00000110, // Color (7, 5, 3) (10, 0)
        8'b00110100, // Color (9, 7, 4) (11, 0)
        8'b00110010, // Color (4, 3, 2) (12, 0)
        8'b00110100, // Color (9, 7, 4) (13, 0)
        8'b00000110, // Color (7, 5, 3) (14, 0)
        8'b00111000, // Color (5, 4, 2) (15, 0)
        8'b00000110, // Color (7, 5, 3) (0, 1)
        8'b00110010, // Color (4, 3, 2) (1, 1)
        8'b00110100, // Color (9, 7, 4) (2, 1)
        8'b00111000, // Color (5, 4, 2) (3, 1)
        8'b00000110, // Color (7, 5, 3) (4, 1)
        8'b00110110, // Color (3, 2, 1) (5, 1)
        8'b00110100, // Color (9, 7, 4) (6, 1)
        8'b00111000, // Color (5, 4, 2) (7, 1)
        8'b00000110, // Color (7, 5, 3) (8, 1)
        8'b00110110, // Color (3, 2, 1) (9, 1)
        8'b00000110, // Color (7, 5, 3) (10, 1)
        8'b00110100, // Color (9, 7, 4) (11, 1)
        8'b00110010, // Color (4, 3, 2) (12, 1)
        8'b00000110, // Color (7, 5, 3) (13, 1)
        8'b00000110, // Color (7, 5, 3) (14, 1)
        8'b00111000, // Color (5, 4, 2) (15, 1)
        8'b00000110, // Color (7, 5, 3) (0, 2)
        8'b00110110, // Color (3, 2, 1) (1, 2)
        8'b00111000, // Color (5, 4, 2) (2, 2)
        8'b00111000, // Color (5, 4, 2) (3, 2)
        8'b00000110, // Color (7, 5, 3) (4, 2)
        8'b00110110, // Color (3, 2, 1) (5, 2)
        8'b00110100, // Color (9, 7, 4) (6, 2)
        8'b00111000, // Color (5, 4, 2) (7, 2)
        8'b00000110, // Color (7, 5, 3) (8, 2)
        8'b00110010, // Color (4, 3, 2) (9, 2)
        8'b00000110, // Color (7, 5, 3) (10, 2)
        8'b00110010, // Color (4, 3, 2) (11, 2)
        8'b00110010, // Color (4, 3, 2) (12, 2)
        8'b00000110, // Color (7, 5, 3) (13, 2)
        8'b00000110, // Color (7, 5, 3) (14, 2)
        8'b00111000, // Color (5, 4, 2) (15, 2)
        8'b00110100, // Color (9, 7, 4) (0, 3)
        8'b00110110, // Color (3, 2, 1) (1, 3)
        8'b00000110, // Color (7, 5, 3) (2, 3)
        8'b00111000, // Color (5, 4, 2) (3, 3)
        8'b00000110, // Color (7, 5, 3) (4, 3)
        8'b00110010, // Color (4, 3, 2) (5, 3)
        8'b00000110, // Color (7, 5, 3) (6, 3)
        8'b00111000, // Color (5, 4, 2) (7, 3)
        8'b00000110, // Color (7, 5, 3) (8, 3)
        8'b00111000, // Color (5, 4, 2) (9, 3)
        8'b00000110, // Color (7, 5, 3) (10, 3)
        8'b00110110, // Color (3, 2, 1) (11, 3)
        8'b00110010, // Color (4, 3, 2) (12, 3)
        8'b00000110, // Color (7, 5, 3) (13, 3)
        8'b00110100, // Color (9, 7, 4) (14, 3)
        8'b00111000, // Color (5, 4, 2) (15, 3)
        8'b00110100, // Color (9, 7, 4) (0, 4)
        8'b00110010, // Color (4, 3, 2) (1, 4)
        8'b00000110, // Color (7, 5, 3) (2, 4)
        8'b00111000, // Color (5, 4, 2) (3, 4)
        8'b00000110, // Color (7, 5, 3) (4, 4)
        8'b00110110, // Color (3, 2, 1) (5, 4)
        8'b00000110, // Color (7, 5, 3) (6, 4)
        8'b00111000, // Color (5, 4, 2) (7, 4)
        8'b00110100, // Color (9, 7, 4) (8, 4)
        8'b00111000, // Color (5, 4, 2) (9, 4)
        8'b00000110, // Color (7, 5, 3) (10, 4)
        8'b00111000, // Color (5, 4, 2) (11, 4)
        8'b00000110, // Color (7, 5, 3) (12, 4)
        8'b00110010, // Color (4, 3, 2) (13, 4)
        8'b00110100, // Color (9, 7, 4) (14, 4)
        8'b00000110, // Color (7, 5, 3) (15, 4)
        8'b00110100, // Color (9, 7, 4) (0, 5)
        8'b00000110, // Color (7, 5, 3) (1, 5)
        8'b00110010, // Color (4, 3, 2) (2, 5)
        8'b00000110, // Color (7, 5, 3) (3, 5)
        8'b00110100, // Color (9, 7, 4) (4, 5)
        8'b00110010, // Color (4, 3, 2) (5, 5)
        8'b00000110, // Color (7, 5, 3) (6, 5)
        8'b00110010, // Color (4, 3, 2) (7, 5)
        8'b00110100, // Color (9, 7, 4) (8, 5)
        8'b00111000, // Color (5, 4, 2) (9, 5)
        8'b00110100, // Color (9, 7, 4) (10, 5)
        8'b00110010, // Color (4, 3, 2) (11, 5)
        8'b00000110, // Color (7, 5, 3) (12, 5)
        8'b00110010, // Color (4, 3, 2) (13, 5)
        8'b00110100, // Color (9, 7, 4) (14, 5)
        8'b00000110, // Color (7, 5, 3) (15, 5)
        8'b00111000, // Color (5, 4, 2) (0, 6)
        8'b00000110, // Color (7, 5, 3) (1, 6)
        8'b00110010, // Color (4, 3, 2) (2, 6)
        8'b00000110, // Color (7, 5, 3) (3, 6)
        8'b00110100, // Color (9, 7, 4) (4, 6)
        8'b00111000, // Color (5, 4, 2) (5, 6)
        8'b00111000, // Color (5, 4, 2) (6, 6)
        8'b00000110, // Color (7, 5, 3) (7, 6)
        8'b00110100, // Color (9, 7, 4) (8, 6)
        8'b00000110, // Color (7, 5, 3) (9, 6)
        8'b00110100, // Color (9, 7, 4) (10, 6)
        8'b00000110, // Color (7, 5, 3) (11, 6)
        8'b00000110, // Color (7, 5, 3) (12, 6)
        8'b00110010, // Color (4, 3, 2) (13, 6)
        8'b00110100, // Color (9, 7, 4) (14, 6)
        8'b00000110, // Color (7, 5, 3) (15, 6)
        8'b00111000, // Color (5, 4, 2) (0, 7)
        8'b00000110, // Color (7, 5, 3) (1, 7)
        8'b00110110, // Color (3, 2, 1) (2, 7)
        8'b00000110, // Color (7, 5, 3) (3, 7)
        8'b00110100, // Color (9, 7, 4) (4, 7)
        8'b00000110, // Color (7, 5, 3) (5, 7)
        8'b00111000, // Color (5, 4, 2) (6, 7)
        8'b00110100, // Color (9, 7, 4) (7, 7)
        8'b00000110, // Color (7, 5, 3) (8, 7)
        8'b00000110, // Color (7, 5, 3) (9, 7)
        8'b00110100, // Color (9, 7, 4) (10, 7)
        8'b00111000, // Color (5, 4, 2) (11, 7)
        8'b00000110, // Color (7, 5, 3) (12, 7)
        8'b00111000, // Color (5, 4, 2) (13, 7)
        8'b00110100, // Color (9, 7, 4) (14, 7)
        8'b00000110, // Color (7, 5, 3) (15, 7)
        8'b00000110, // Color (7, 5, 3) (0, 8)
        8'b00110010, // Color (4, 3, 2) (1, 8)
        8'b00110110, // Color (3, 2, 1) (2, 8)
        8'b00110100, // Color (9, 7, 4) (3, 8)
        8'b00000110, // Color (7, 5, 3) (4, 8)
        8'b00000110, // Color (7, 5, 3) (5, 8)
        8'b00111000, // Color (5, 4, 2) (6, 8)
        8'b00110100, // Color (9, 7, 4) (7, 8)
        8'b00000110, // Color (7, 5, 3) (8, 8)
        8'b00111000, // Color (5, 4, 2) (9, 8)
        8'b00110100, // Color (9, 7, 4) (10, 8)
        8'b00111000, // Color (5, 4, 2) (11, 8)
        8'b00110100, // Color (9, 7, 4) (12, 8)
        8'b00111000, // Color (5, 4, 2) (13, 8)
        8'b00110100, // Color (9, 7, 4) (14, 8)
        8'b00000110, // Color (7, 5, 3) (15, 8)
        8'b00000110, // Color (7, 5, 3) (0, 9)
        8'b00000110, // Color (7, 5, 3) (1, 9)
        8'b00110010, // Color (4, 3, 2) (2, 9)
        8'b00110100, // Color (9, 7, 4) (3, 9)
        8'b00000110, // Color (7, 5, 3) (4, 9)
        8'b00000110, // Color (7, 5, 3) (5, 9)
        8'b00111000, // Color (5, 4, 2) (6, 9)
        8'b00000110, // Color (7, 5, 3) (7, 9)
        8'b00000110, // Color (7, 5, 3) (8, 9)
        8'b00111000, // Color (5, 4, 2) (9, 9)
        8'b00110100, // Color (9, 7, 4) (10, 9)
        8'b00110010, // Color (4, 3, 2) (11, 9)
        8'b00110100, // Color (9, 7, 4) (12, 9)
        8'b00000110, // Color (7, 5, 3) (13, 9)
        8'b00110110, // Color (3, 2, 1) (14, 9)
        8'b00000110, // Color (7, 5, 3) (15, 9)
        8'b00000110, // Color (7, 5, 3) (0, 10)
        8'b00000110, // Color (7, 5, 3) (1, 10)
        8'b00000110, // Color (7, 5, 3) (2, 10)
        8'b00110100, // Color (9, 7, 4) (3, 10)
        8'b00000110, // Color (7, 5, 3) (4, 10)
        8'b00111000, // Color (5, 4, 2) (5, 10)
        8'b00000110, // Color (7, 5, 3) (6, 10)
        8'b00110110, // Color (3, 2, 1) (7, 10)
        8'b00000110, // Color (7, 5, 3) (8, 10)
        8'b00111000, // Color (5, 4, 2) (9, 10)
        8'b00000110, // Color (7, 5, 3) (10, 10)
        8'b00110010, // Color (4, 3, 2) (11, 10)
        8'b00110100, // Color (9, 7, 4) (12, 10)
        8'b00000110, // Color (7, 5, 3) (13, 10)
        8'b00110110, // Color (3, 2, 1) (14, 10)
        8'b00000110, // Color (7, 5, 3) (15, 10)
        8'b00000110, // Color (7, 5, 3) (0, 11)
        8'b00110010, // Color (4, 3, 2) (1, 11)
        8'b00000110, // Color (7, 5, 3) (2, 11)
        8'b00110100, // Color (9, 7, 4) (3, 11)
        8'b00000110, // Color (7, 5, 3) (4, 11)
        8'b00111000, // Color (5, 4, 2) (5, 11)
        8'b00000110, // Color (7, 5, 3) (6, 11)
        8'b00110110, // Color (3, 2, 1) (7, 11)
        8'b00110100, // Color (9, 7, 4) (8, 11)
        8'b00000110, // Color (7, 5, 3) (9, 11)
        8'b00000110, // Color (7, 5, 3) (10, 11)
        8'b00110110, // Color (3, 2, 1) (11, 11)
        8'b00110100, // Color (9, 7, 4) (12, 11)
        8'b00000110, // Color (7, 5, 3) (13, 11)
        8'b00110010, // Color (4, 3, 2) (14, 11)
        8'b00000110, // Color (7, 5, 3) (15, 11)
        8'b00110100, // Color (9, 7, 4) (0, 12)
        8'b00110010, // Color (4, 3, 2) (1, 12)
        8'b00000110, // Color (7, 5, 3) (2, 12)
        8'b00000110, // Color (7, 5, 3) (3, 12)
        8'b00110100, // Color (9, 7, 4) (4, 12)
        8'b00111000, // Color (5, 4, 2) (5, 12)
        8'b00110100, // Color (9, 7, 4) (6, 12)
        8'b00110110, // Color (3, 2, 1) (7, 12)
        8'b00110100, // Color (9, 7, 4) (8, 12)
        8'b00111000, // Color (5, 4, 2) (9, 12)
        8'b00000110, // Color (7, 5, 3) (10, 12)
        8'b00110110, // Color (3, 2, 1) (11, 12)
        8'b00000110, // Color (7, 5, 3) (12, 12)
        8'b00000110, // Color (7, 5, 3) (13, 12)
        8'b00111000, // Color (5, 4, 2) (14, 12)
        8'b00000110, // Color (7, 5, 3) (15, 12)
        8'b00110100, // Color (9, 7, 4) (0, 13)
        8'b00000110, // Color (7, 5, 3) (1, 13)
        8'b00110010, // Color (4, 3, 2) (2, 13)
        8'b00000110, // Color (7, 5, 3) (3, 13)
        8'b00110100, // Color (9, 7, 4) (4, 13)
        8'b00000110, // Color (7, 5, 3) (5, 13)
        8'b00000110, // Color (7, 5, 3) (6, 13)
        8'b00110010, // Color (4, 3, 2) (7, 13)
        8'b00110100, // Color (9, 7, 4) (8, 13)
        8'b00111000, // Color (5, 4, 2) (9, 13)
        8'b00000110, // Color (7, 5, 3) (10, 13)
        8'b00110010, // Color (4, 3, 2) (11, 13)
        8'b00000110, // Color (7, 5, 3) (12, 13)
        8'b00000110, // Color (7, 5, 3) (13, 13)
        8'b00000110, // Color (7, 5, 3) (14, 13)
        8'b00000110, // Color (7, 5, 3) (15, 13)
        8'b00110100, // Color (9, 7, 4) (0, 14)
        8'b00000110, // Color (7, 5, 3) (1, 14)
        8'b00110010, // Color (4, 3, 2) (2, 14)
        8'b00110100, // Color (9, 7, 4) (3, 14)
        8'b00000110, // Color (7, 5, 3) (4, 14)
        8'b00000110, // Color (7, 5, 3) (5, 14)
        8'b00110100, // Color (9, 7, 4) (6, 14)
        8'b00110110, // Color (3, 2, 1) (7, 14)
        8'b00000110, // Color (7, 5, 3) (8, 14)
        8'b00110010, // Color (4, 3, 2) (9, 14)
        8'b00000110, // Color (7, 5, 3) (10, 14)
        8'b00110010, // Color (4, 3, 2) (11, 14)
        8'b00110010, // Color (4, 3, 2) (12, 14)
        8'b00110100, // Color (9, 7, 4) (13, 14)
        8'b00000110, // Color (7, 5, 3) (14, 14)
        8'b00000110, // Color (7, 5, 3) (15, 14)
        8'b00110100, // Color (9, 7, 4) (0, 15)
        8'b00000110, // Color (7, 5, 3) (1, 15)
        8'b00110010, // Color (4, 3, 2) (2, 15)
        8'b00110100, // Color (9, 7, 4) (3, 15)
        8'b00110010, // Color (4, 3, 2) (4, 15)
        8'b00000110, // Color (7, 5, 3) (5, 15)
        8'b00110100, // Color (9, 7, 4) (6, 15)
        8'b00110010, // Color (4, 3, 2) (7, 15)
        8'b00000110, // Color (7, 5, 3) (8, 15)
        8'b00110010, // Color (4, 3, 2) (9, 15)
        8'b00000110, // Color (7, 5, 3) (10, 15)
        8'b00000110, // Color (7, 5, 3) (11, 15)
        8'b00110010, // Color (4, 3, 2) (12, 15)
        8'b00110100, // Color (9, 7, 4) (13, 15)
        8'b00000110, // Color (7, 5, 3) (14, 15)
        8'b00111000, // Color (5, 4, 2) (15, 15)
        // 04_oak_log_top
        8'b00111000, // Color (5, 4, 2) (0, 0)
        8'b00110010, // Color (4, 3, 2) (1, 0)
        8'b00111000, // Color (5, 4, 2) (2, 0)
        8'b00000110, // Color (7, 5, 3) (3, 0)
        8'b00111000, // Color (5, 4, 2) (4, 0)
        8'b00110010, // Color (4, 3, 2) (5, 0)
        8'b00111000, // Color (5, 4, 2) (6, 0)
        8'b00111000, // Color (5, 4, 2) (7, 0)
        8'b00000110, // Color (7, 5, 3) (8, 0)
        8'b00110010, // Color (4, 3, 2) (9, 0)
        8'b00111000, // Color (5, 4, 2) (10, 0)
        8'b00111000, // Color (5, 4, 2) (11, 0)
        8'b00110010, // Color (4, 3, 2) (12, 0)
        8'b00111000, // Color (5, 4, 2) (13, 0)
        8'b00111000, // Color (5, 4, 2) (14, 0)
        8'b00111000, // Color (5, 4, 2) (15, 0)
        8'b00110010, // Color (4, 3, 2) (0, 1)
        8'b00111010, // Color (11, 9, 5) (1, 1)
        8'b00111010, // Color (11, 9, 5) (2, 1)
        8'b00111010, // Color (11, 9, 5) (3, 1)
        8'b00111010, // Color (11, 9, 5) (4, 1)
        8'b00111100, // Color (10, 8, 5) (5, 1)
        8'b00111010, // Color (11, 9, 5) (6, 1)
        8'b00111100, // Color (10, 8, 5) (7, 1)
        8'b00111110, // Color (12, 9, 6) (8, 1)
        8'b00111100, // Color (10, 8, 5) (9, 1)
        8'b00111100, // Color (10, 8, 5) (10, 1)
        8'b00111010, // Color (11, 9, 5) (11, 1)
        8'b00111010, // Color (11, 9, 5) (12, 1)
        8'b00111010, // Color (11, 9, 5) (13, 1)
        8'b00111010, // Color (11, 9, 5) (14, 1)
        8'b00110010, // Color (4, 3, 2) (15, 1)
        8'b00111000, // Color (5, 4, 2) (0, 2)
        8'b00111010, // Color (11, 9, 5) (1, 2)
        8'b01000000, // Color (7, 6, 3) (2, 2)
        8'b01000000, // Color (7, 6, 3) (3, 2)
        8'b00110100, // Color (9, 7, 4) (4, 2)
        8'b00110100, // Color (9, 7, 4) (5, 2)
        8'b01000010, // Color (9, 8, 4) (6, 2)
        8'b00110100, // Color (9, 7, 4) (7, 2)
        8'b01000010, // Color (9, 8, 4) (8, 2)
        8'b01000010, // Color (9, 8, 4) (9, 2)
        8'b01000010, // Color (9, 8, 4) (10, 2)
        8'b01000010, // Color (9, 8, 4) (11, 2)
        8'b00110100, // Color (9, 7, 4) (12, 2)
        8'b00110100, // Color (9, 7, 4) (13, 2)
        8'b00111110, // Color (12, 9, 6) (14, 2)
        8'b00111000, // Color (5, 4, 2) (15, 2)
        8'b00111000, // Color (5, 4, 2) (0, 3)
        8'b00111010, // Color (11, 9, 5) (1, 3)
        8'b01000000, // Color (7, 6, 3) (2, 3)
        8'b00111110, // Color (12, 9, 6) (3, 3)
        8'b00111110, // Color (12, 9, 6) (4, 3)
        8'b00111010, // Color (11, 9, 5) (5, 3)
        8'b00111010, // Color (11, 9, 5) (6, 3)
        8'b00111010, // Color (11, 9, 5) (7, 3)
        8'b00111010, // Color (11, 9, 5) (8, 3)
        8'b00111100, // Color (10, 8, 5) (9, 3)
        8'b00111010, // Color (11, 9, 5) (10, 3)
        8'b00111010, // Color (11, 9, 5) (11, 3)
        8'b00111010, // Color (11, 9, 5) (12, 3)
        8'b00110100, // Color (9, 7, 4) (13, 3)
        8'b00111010, // Color (11, 9, 5) (14, 3)
        8'b00111000, // Color (5, 4, 2) (15, 3)
        8'b00111000, // Color (5, 4, 2) (0, 4)
        8'b00111100, // Color (10, 8, 5) (1, 4)
        8'b00110100, // Color (9, 7, 4) (2, 4)
        8'b00111010, // Color (11, 9, 5) (3, 4)
        8'b00111100, // Color (10, 8, 5) (4, 4)
        8'b00111100, // Color (10, 8, 5) (5, 4)
        8'b00111100, // Color (10, 8, 5) (6, 4)
        8'b00111100, // Color (10, 8, 5) (7, 4)
        8'b00111100, // Color (10, 8, 5) (8, 4)
        8'b00111100, // Color (10, 8, 5) (9, 4)
        8'b00111100, // Color (10, 8, 5) (10, 4)
        8'b00111100, // Color (10, 8, 5) (11, 4)
        8'b00111010, // Color (11, 9, 5) (12, 4)
        8'b01000010, // Color (9, 8, 4) (13, 4)
        8'b00111100, // Color (10, 8, 5) (14, 4)
        8'b00111000, // Color (5, 4, 2) (15, 4)
        8'b00110010, // Color (4, 3, 2) (0, 5)
        8'b00111010, // Color (11, 9, 5) (1, 5)
        8'b01000010, // Color (9, 8, 4) (2, 5)
        8'b00111010, // Color (11, 9, 5) (3, 5)
        8'b00111100, // Color (10, 8, 5) (4, 5)
        8'b00110100, // Color (9, 7, 4) (5, 5)
        8'b00110100, // Color (9, 7, 4) (6, 5)
        8'b01000010, // Color (9, 8, 4) (7, 5)
        8'b01000010, // Color (9, 8, 4) (8, 5)
        8'b00110100, // Color (9, 7, 4) (9, 5)
        8'b00110100, // Color (9, 7, 4) (10, 5)
        8'b00111100, // Color (10, 8, 5) (11, 5)
        8'b00111010, // Color (11, 9, 5) (12, 5)
        8'b00110100, // Color (9, 7, 4) (13, 5)
        8'b00111100, // Color (10, 8, 5) (14, 5)
        8'b00110010, // Color (4, 3, 2) (15, 5)
        8'b00111000, // Color (5, 4, 2) (0, 6)
        8'b00111100, // Color (10, 8, 5) (1, 6)
        8'b00110100, // Color (9, 7, 4) (2, 6)
        8'b00111100, // Color (10, 8, 5) (3, 6)
        8'b00111100, // Color (10, 8, 5) (4, 6)
        8'b01000000, // Color (7, 6, 3) (5, 6)
        8'b00111100, // Color (10, 8, 5) (6, 6)
        8'b00111100, // Color (10, 8, 5) (7, 6)
        8'b00111100, // Color (10, 8, 5) (8, 6)
        8'b00111100, // Color (10, 8, 5) (9, 6)
        8'b00110100, // Color (9, 7, 4) (10, 6)
        8'b00111100, // Color (10, 8, 5) (11, 6)
        8'b00111100, // Color (10, 8, 5) (12, 6)
        8'b00110100, // Color (9, 7, 4) (13, 6)
        8'b00111010, // Color (11, 9, 5) (14, 6)
        8'b00111000, // Color (5, 4, 2) (15, 6)
        8'b00111000, // Color (5, 4, 2) (0, 7)
        8'b00111100, // Color (10, 8, 5) (1, 7)
        8'b01000010, // Color (9, 8, 4) (2, 7)
        8'b00111010, // Color (11, 9, 5) (3, 7)
        8'b00111100, // Color (10, 8, 5) (4, 7)
        8'b00110100, // Color (9, 7, 4) (5, 7)
        8'b00111100, // Color (10, 8, 5) (6, 7)
        8'b01000010, // Color (9, 8, 4) (7, 7)
        8'b01000010, // Color (9, 8, 4) (8, 7)
        8'b00111100, // Color (10, 8, 5) (9, 7)
        8'b01000010, // Color (9, 8, 4) (10, 7)
        8'b00111100, // Color (10, 8, 5) (11, 7)
        8'b00111010, // Color (11, 9, 5) (12, 7)
        8'b01000010, // Color (9, 8, 4) (13, 7)
        8'b00111100, // Color (10, 8, 5) (14, 7)
        8'b00111000, // Color (5, 4, 2) (15, 7)
        8'b00111000, // Color (5, 4, 2) (0, 8)
        8'b00111100, // Color (10, 8, 5) (1, 8)
        8'b01000010, // Color (9, 8, 4) (2, 8)
        8'b00111010, // Color (11, 9, 5) (3, 8)
        8'b00111100, // Color (10, 8, 5) (4, 8)
        8'b00110100, // Color (9, 7, 4) (5, 8)
        8'b00111100, // Color (10, 8, 5) (6, 8)
        8'b01000010, // Color (9, 8, 4) (7, 8)
        8'b00110100, // Color (9, 7, 4) (8, 8)
        8'b00111100, // Color (10, 8, 5) (9, 8)
        8'b00110100, // Color (9, 7, 4) (10, 8)
        8'b00111100, // Color (10, 8, 5) (11, 8)
        8'b00111010, // Color (11, 9, 5) (12, 8)
        8'b00110100, // Color (9, 7, 4) (13, 8)
        8'b00111100, // Color (10, 8, 5) (14, 8)
        8'b00111000, // Color (5, 4, 2) (15, 8)
        8'b00110010, // Color (4, 3, 2) (0, 9)
        8'b00111100, // Color (10, 8, 5) (1, 9)
        8'b01000010, // Color (9, 8, 4) (2, 9)
        8'b00111010, // Color (11, 9, 5) (3, 9)
        8'b00111100, // Color (10, 8, 5) (4, 9)
        8'b00110100, // Color (9, 7, 4) (5, 9)
        8'b00111100, // Color (10, 8, 5) (6, 9)
        8'b00111100, // Color (10, 8, 5) (7, 9)
        8'b00111100, // Color (10, 8, 5) (8, 9)
        8'b00111100, // Color (10, 8, 5) (9, 9)
        8'b01000010, // Color (9, 8, 4) (10, 9)
        8'b00111100, // Color (10, 8, 5) (11, 9)
        8'b00111100, // Color (10, 8, 5) (12, 9)
        8'b00110100, // Color (9, 7, 4) (13, 9)
        8'b00111100, // Color (10, 8, 5) (14, 9)
        8'b00110010, // Color (4, 3, 2) (15, 9)
        8'b00111000, // Color (5, 4, 2) (0, 10)
        8'b00111100, // Color (10, 8, 5) (1, 10)
        8'b00110100, // Color (9, 7, 4) (2, 10)
        8'b00111010, // Color (11, 9, 5) (3, 10)
        8'b00111100, // Color (10, 8, 5) (4, 10)
        8'b00110100, // Color (9, 7, 4) (5, 10)
        8'b00110100, // Color (9, 7, 4) (6, 10)
        8'b01000000, // Color (7, 6, 3) (7, 10)
        8'b00110100, // Color (9, 7, 4) (8, 10)
        8'b01000010, // Color (9, 8, 4) (9, 10)
        8'b01000010, // Color (9, 8, 4) (10, 10)
        8'b00111100, // Color (10, 8, 5) (11, 10)
        8'b00111010, // Color (11, 9, 5) (12, 10)
        8'b01000010, // Color (9, 8, 4) (13, 10)
        8'b00111100, // Color (10, 8, 5) (14, 10)
        8'b00111000, // Color (5, 4, 2) (15, 10)
        8'b00111000, // Color (5, 4, 2) (0, 11)
        8'b00111100, // Color (10, 8, 5) (1, 11)
        8'b01000010, // Color (9, 8, 4) (2, 11)
        8'b00111010, // Color (11, 9, 5) (3, 11)
        8'b00111100, // Color (10, 8, 5) (4, 11)
        8'b00111100, // Color (10, 8, 5) (5, 11)
        8'b00111100, // Color (10, 8, 5) (6, 11)
        8'b00111100, // Color (10, 8, 5) (7, 11)
        8'b00111100, // Color (10, 8, 5) (8, 11)
        8'b00111100, // Color (10, 8, 5) (9, 11)
        8'b00111100, // Color (10, 8, 5) (10, 11)
        8'b00111100, // Color (10, 8, 5) (11, 11)
        8'b00111010, // Color (11, 9, 5) (12, 11)
        8'b00110100, // Color (9, 7, 4) (13, 11)
        8'b00111100, // Color (10, 8, 5) (14, 11)
        8'b00111000, // Color (5, 4, 2) (15, 11)
        8'b00110010, // Color (4, 3, 2) (0, 12)
        8'b00111010, // Color (11, 9, 5) (1, 12)
        8'b01000010, // Color (9, 8, 4) (2, 12)
        8'b00111010, // Color (11, 9, 5) (3, 12)
        8'b00111010, // Color (11, 9, 5) (4, 12)
        8'b00111100, // Color (10, 8, 5) (5, 12)
        8'b00111010, // Color (11, 9, 5) (6, 12)
        8'b00111010, // Color (11, 9, 5) (7, 12)
        8'b00111010, // Color (11, 9, 5) (8, 12)
        8'b00111010, // Color (11, 9, 5) (9, 12)
        8'b00111010, // Color (11, 9, 5) (10, 12)
        8'b00111110, // Color (12, 9, 6) (11, 12)
        8'b00111010, // Color (11, 9, 5) (12, 12)
        8'b00110100, // Color (9, 7, 4) (13, 12)
        8'b00111100, // Color (10, 8, 5) (14, 12)
        8'b00110010, // Color (4, 3, 2) (15, 12)
        8'b00111000, // Color (5, 4, 2) (0, 13)
        8'b00111010, // Color (11, 9, 5) (1, 13)
        8'b01000010, // Color (9, 8, 4) (2, 13)
        8'b00110100, // Color (9, 7, 4) (3, 13)
        8'b01000010, // Color (9, 8, 4) (4, 13)
        8'b00110100, // Color (9, 7, 4) (5, 13)
        8'b00110100, // Color (9, 7, 4) (6, 13)
        8'b00110100, // Color (9, 7, 4) (7, 13)
        8'b00110100, // Color (9, 7, 4) (8, 13)
        8'b00110100, // Color (9, 7, 4) (9, 13)
        8'b00110100, // Color (9, 7, 4) (10, 13)
        8'b00110100, // Color (9, 7, 4) (11, 13)
        8'b00110100, // Color (9, 7, 4) (12, 13)
        8'b00110100, // Color (9, 7, 4) (13, 13)
        8'b00111010, // Color (11, 9, 5) (14, 13)
        8'b00111000, // Color (5, 4, 2) (15, 13)
        8'b00111000, // Color (5, 4, 2) (0, 14)
        8'b00111010, // Color (11, 9, 5) (1, 14)
        8'b00111010, // Color (11, 9, 5) (2, 14)
        8'b00111010, // Color (11, 9, 5) (3, 14)
        8'b00111100, // Color (10, 8, 5) (4, 14)
        8'b00111100, // Color (10, 8, 5) (5, 14)
        8'b00111010, // Color (11, 9, 5) (6, 14)
        8'b00111100, // Color (10, 8, 5) (7, 14)
        8'b00111100, // Color (10, 8, 5) (8, 14)
        8'b00111110, // Color (12, 9, 6) (9, 14)
        8'b00111100, // Color (10, 8, 5) (10, 14)
        8'b00111100, // Color (10, 8, 5) (11, 14)
        8'b00111010, // Color (11, 9, 5) (12, 14)
        8'b00111010, // Color (11, 9, 5) (13, 14)
        8'b00111010, // Color (11, 9, 5) (14, 14)
        8'b00111000, // Color (5, 4, 2) (15, 14)
        8'b00111000, // Color (5, 4, 2) (0, 15)
        8'b00110010, // Color (4, 3, 2) (1, 15)
        8'b00111000, // Color (5, 4, 2) (2, 15)
        8'b00111000, // Color (5, 4, 2) (3, 15)
        8'b00111000, // Color (5, 4, 2) (4, 15)
        8'b00110010, // Color (4, 3, 2) (5, 15)
        8'b00111000, // Color (5, 4, 2) (6, 15)
        8'b00111000, // Color (5, 4, 2) (7, 15)
        8'b00000110, // Color (7, 5, 3) (8, 15)
        8'b00110010, // Color (4, 3, 2) (9, 15)
        8'b00111000, // Color (5, 4, 2) (10, 15)
        8'b00111000, // Color (5, 4, 2) (11, 15)
        8'b00110010, // Color (4, 3, 2) (12, 15)
        8'b00000110, // Color (7, 5, 3) (13, 15)
        8'b00111000, // Color (5, 4, 2) (14, 15)
        8'b00111000, // Color (5, 4, 2) (15, 15)
        // 05_oak_planks
        8'b00111010, // Color (11, 9, 5) (0, 0)
        8'b00111100, // Color (10, 8, 5) (1, 0)
        8'b00111010, // Color (11, 9, 5) (2, 0)
        8'b00111110, // Color (12, 9, 6) (3, 0)
        8'b00111110, // Color (12, 9, 6) (4, 0)
        8'b00111110, // Color (12, 9, 6) (5, 0)
        8'b00111110, // Color (12, 9, 6) (6, 0)
        8'b00111110, // Color (12, 9, 6) (7, 0)
        8'b00111010, // Color (11, 9, 5) (8, 0)
        8'b00111110, // Color (12, 9, 6) (9, 0)
        8'b00111110, // Color (12, 9, 6) (10, 0)
        8'b00111110, // Color (12, 9, 6) (11, 0)
        8'b00111110, // Color (12, 9, 6) (12, 0)
        8'b00111110, // Color (12, 9, 6) (13, 0)
        8'b00111010, // Color (11, 9, 5) (14, 0)
        8'b00110100, // Color (9, 7, 4) (15, 0)
        8'b00111010, // Color (11, 9, 5) (0, 1)
        8'b00111010, // Color (11, 9, 5) (1, 1)
        8'b00111100, // Color (10, 8, 5) (2, 1)
        8'b00111100, // Color (10, 8, 5) (3, 1)
        8'b00110100, // Color (9, 7, 4) (4, 1)
        8'b01000010, // Color (9, 8, 4) (5, 1)
        8'b00111100, // Color (10, 8, 5) (6, 1)
        8'b00111010, // Color (11, 9, 5) (7, 1)
        8'b00111010, // Color (11, 9, 5) (8, 1)
        8'b00111010, // Color (11, 9, 5) (9, 1)
        8'b00111100, // Color (10, 8, 5) (10, 1)
        8'b00111100, // Color (10, 8, 5) (11, 1)
        8'b00111010, // Color (11, 9, 5) (12, 1)
        8'b00111010, // Color (11, 9, 5) (13, 1)
        8'b01000010, // Color (9, 8, 4) (14, 1)
        8'b01000010, // Color (9, 8, 4) (15, 1)
        8'b00111100, // Color (10, 8, 5) (0, 2)
        8'b00111010, // Color (11, 9, 5) (1, 2)
        8'b00111010, // Color (11, 9, 5) (2, 2)
        8'b00111010, // Color (11, 9, 5) (3, 2)
        8'b00111100, // Color (10, 8, 5) (4, 2)
        8'b00111010, // Color (11, 9, 5) (5, 2)
        8'b00111100, // Color (10, 8, 5) (6, 2)
        8'b01000010, // Color (9, 8, 4) (7, 2)
        8'b01000010, // Color (9, 8, 4) (8, 2)
        8'b01000010, // Color (9, 8, 4) (9, 2)
        8'b01000010, // Color (9, 8, 4) (10, 2)
        8'b00111100, // Color (10, 8, 5) (11, 2)
        8'b00111100, // Color (10, 8, 5) (12, 2)
        8'b00111010, // Color (11, 9, 5) (13, 2)
        8'b00111010, // Color (11, 9, 5) (14, 2)
        8'b00110100, // Color (9, 7, 4) (15, 2)
        8'b00110100, // Color (9, 7, 4) (0, 3)
        8'b01000000, // Color (7, 6, 3) (1, 3)
        8'b01000000, // Color (7, 6, 3) (2, 3)
        8'b00110100, // Color (9, 7, 4) (3, 3)
        8'b00110100, // Color (9, 7, 4) (4, 3)
        8'b01000000, // Color (7, 6, 3) (5, 3)
        8'b01000100, // Color (6, 5, 2) (6, 3)
        8'b01000100, // Color (6, 5, 2) (7, 3)
        8'b01000000, // Color (7, 6, 3) (8, 3)
        8'b01000000, // Color (7, 6, 3) (9, 3)
        8'b01000100, // Color (6, 5, 2) (10, 3)
        8'b01000000, // Color (7, 6, 3) (11, 3)
        8'b01000100, // Color (6, 5, 2) (12, 3)
        8'b01000100, // Color (6, 5, 2) (13, 3)
        8'b01000000, // Color (7, 6, 3) (14, 3)
        8'b01000100, // Color (6, 5, 2) (15, 3)
        8'b00111010, // Color (11, 9, 5) (0, 4)
        8'b00111110, // Color (12, 9, 6) (1, 4)
        8'b01000010, // Color (9, 8, 4) (2, 4)
        8'b00111110, // Color (12, 9, 6) (3, 4)
        8'b00111110, // Color (12, 9, 6) (4, 4)
        8'b00111110, // Color (12, 9, 6) (5, 4)
        8'b00111110, // Color (12, 9, 6) (6, 4)
        8'b01000010, // Color (9, 8, 4) (7, 4)
        8'b00111110, // Color (12, 9, 6) (8, 4)
        8'b00111110, // Color (12, 9, 6) (9, 4)
        8'b00111110, // Color (12, 9, 6) (10, 4)
        8'b00111010, // Color (11, 9, 5) (11, 4)
        8'b00111100, // Color (10, 8, 5) (12, 4)
        8'b00111100, // Color (10, 8, 5) (13, 4)
        8'b01000010, // Color (9, 8, 4) (14, 4)
        8'b00111010, // Color (11, 9, 5) (15, 4)
        8'b00111100, // Color (10, 8, 5) (0, 5)
        8'b00111010, // Color (11, 9, 5) (1, 5)
        8'b00111010, // Color (11, 9, 5) (2, 5)
        8'b00111100, // Color (10, 8, 5) (3, 5)
        8'b01000010, // Color (9, 8, 4) (4, 5)
        8'b00111100, // Color (10, 8, 5) (5, 5)
        8'b01000010, // Color (9, 8, 4) (6, 5)
        8'b00110100, // Color (9, 7, 4) (7, 5)
        8'b01000010, // Color (9, 8, 4) (8, 5)
        8'b00111100, // Color (10, 8, 5) (9, 5)
        8'b00111100, // Color (10, 8, 5) (10, 5)
        8'b00111010, // Color (11, 9, 5) (11, 5)
        8'b00111010, // Color (11, 9, 5) (12, 5)
        8'b00111010, // Color (11, 9, 5) (13, 5)
        8'b00111010, // Color (11, 9, 5) (14, 5)
        8'b00111100, // Color (10, 8, 5) (15, 5)
        8'b01000010, // Color (9, 8, 4) (0, 6)
        8'b01000010, // Color (9, 8, 4) (1, 6)
        8'b00111100, // Color (10, 8, 5) (2, 6)
        8'b00111010, // Color (11, 9, 5) (3, 6)
        8'b00111100, // Color (10, 8, 5) (4, 6)
        8'b00111100, // Color (10, 8, 5) (5, 6)
        8'b00111100, // Color (10, 8, 5) (6, 6)
        8'b00110100, // Color (9, 7, 4) (7, 6)
        8'b00111010, // Color (11, 9, 5) (8, 6)
        8'b00111010, // Color (11, 9, 5) (9, 6)
        8'b00111010, // Color (11, 9, 5) (10, 6)
        8'b00111100, // Color (10, 8, 5) (11, 6)
        8'b00111100, // Color (10, 8, 5) (12, 6)
        8'b01000010, // Color (9, 8, 4) (13, 6)
        8'b01000010, // Color (9, 8, 4) (14, 6)
        8'b01000010, // Color (9, 8, 4) (15, 6)
        8'b01000100, // Color (6, 5, 2) (0, 7)
        8'b01000100, // Color (6, 5, 2) (1, 7)
        8'b01000000, // Color (7, 6, 3) (2, 7)
        8'b01000000, // Color (7, 6, 3) (3, 7)
        8'b00110100, // Color (9, 7, 4) (4, 7)
        8'b01000000, // Color (7, 6, 3) (5, 7)
        8'b01000100, // Color (6, 5, 2) (6, 7)
        8'b01000100, // Color (6, 5, 2) (7, 7)
        8'b01000100, // Color (6, 5, 2) (8, 7)
        8'b01000100, // Color (6, 5, 2) (9, 7)
        8'b01000000, // Color (7, 6, 3) (10, 7)
        8'b01000000, // Color (7, 6, 3) (11, 7)
        8'b01000000, // Color (7, 6, 3) (12, 7)
        8'b00110100, // Color (9, 7, 4) (13, 7)
        8'b01000000, // Color (7, 6, 3) (14, 7)
        8'b01000100, // Color (6, 5, 2) (15, 7)
        8'b00111010, // Color (11, 9, 5) (0, 8)
        8'b00111110, // Color (12, 9, 6) (1, 8)
        8'b00111110, // Color (12, 9, 6) (2, 8)
        8'b00111010, // Color (11, 9, 5) (3, 8)
        8'b00111100, // Color (10, 8, 5) (4, 8)
        8'b00111100, // Color (10, 8, 5) (5, 8)
        8'b00111110, // Color (12, 9, 6) (6, 8)
        8'b00111110, // Color (12, 9, 6) (7, 8)
        8'b00111110, // Color (12, 9, 6) (8, 8)
        8'b00111110, // Color (12, 9, 6) (9, 8)
        8'b00111110, // Color (12, 9, 6) (10, 8)
        8'b00111110, // Color (12, 9, 6) (11, 8)
        8'b00111110, // Color (12, 9, 6) (12, 8)
        8'b00111110, // Color (12, 9, 6) (13, 8)
        8'b00111010, // Color (11, 9, 5) (14, 8)
        8'b01000010, // Color (9, 8, 4) (15, 8)
        8'b00111010, // Color (11, 9, 5) (0, 9)
        8'b00111100, // Color (10, 8, 5) (1, 9)
        8'b00111010, // Color (11, 9, 5) (2, 9)
        8'b00111010, // Color (11, 9, 5) (3, 9)
        8'b00111010, // Color (11, 9, 5) (4, 9)
        8'b00111010, // Color (11, 9, 5) (5, 9)
        8'b00111100, // Color (10, 8, 5) (6, 9)
        8'b01000010, // Color (9, 8, 4) (7, 9)
        8'b01000010, // Color (9, 8, 4) (8, 9)
        8'b01000010, // Color (9, 8, 4) (9, 9)
        8'b00111100, // Color (10, 8, 5) (10, 9)
        8'b01000010, // Color (9, 8, 4) (11, 9)
        8'b00111100, // Color (10, 8, 5) (12, 9)
        8'b01000010, // Color (9, 8, 4) (13, 9)
        8'b01000010, // Color (9, 8, 4) (14, 9)
        8'b00110100, // Color (9, 7, 4) (15, 9)
        8'b00111110, // Color (12, 9, 6) (0, 10)
        8'b00111010, // Color (11, 9, 5) (1, 10)
        8'b00111100, // Color (10, 8, 5) (2, 10)
        8'b00111100, // Color (10, 8, 5) (3, 10)
        8'b01000010, // Color (9, 8, 4) (4, 10)
        8'b01000010, // Color (9, 8, 4) (5, 10)
        8'b01000010, // Color (9, 8, 4) (6, 10)
        8'b01000010, // Color (9, 8, 4) (7, 10)
        8'b00111100, // Color (10, 8, 5) (8, 10)
        8'b00111100, // Color (10, 8, 5) (9, 10)
        8'b00111100, // Color (10, 8, 5) (10, 10)
        8'b00111100, // Color (10, 8, 5) (11, 10)
        8'b01000010, // Color (9, 8, 4) (12, 10)
        8'b01000010, // Color (9, 8, 4) (13, 10)
        8'b00111010, // Color (11, 9, 5) (14, 10)
        8'b01000010, // Color (9, 8, 4) (15, 10)
        8'b01000100, // Color (6, 5, 2) (0, 11)
        8'b01000100, // Color (6, 5, 2) (1, 11)
        8'b01000000, // Color (7, 6, 3) (2, 11)
        8'b00110100, // Color (9, 7, 4) (3, 11)
        8'b00110100, // Color (9, 7, 4) (4, 11)
        8'b01000000, // Color (7, 6, 3) (5, 11)
        8'b01000100, // Color (6, 5, 2) (6, 11)
        8'b01000100, // Color (6, 5, 2) (7, 11)
        8'b01000100, // Color (6, 5, 2) (8, 11)
        8'b01000000, // Color (7, 6, 3) (9, 11)
        8'b00110100, // Color (9, 7, 4) (10, 11)
        8'b01000000, // Color (7, 6, 3) (11, 11)
        8'b01000000, // Color (7, 6, 3) (12, 11)
        8'b01000100, // Color (6, 5, 2) (13, 11)
        8'b01000100, // Color (6, 5, 2) (14, 11)
        8'b01000100, // Color (6, 5, 2) (15, 11)
        8'b00111110, // Color (12, 9, 6) (0, 12)
        8'b01000010, // Color (9, 8, 4) (1, 12)
        8'b00111010, // Color (11, 9, 5) (2, 12)
        8'b00111110, // Color (12, 9, 6) (3, 12)
        8'b00111110, // Color (12, 9, 6) (4, 12)
        8'b00111010, // Color (11, 9, 5) (5, 12)
        8'b00111010, // Color (11, 9, 5) (6, 12)
        8'b01000010, // Color (9, 8, 4) (7, 12)
        8'b00111110, // Color (12, 9, 6) (8, 12)
        8'b00111110, // Color (12, 9, 6) (9, 12)
        8'b00111110, // Color (12, 9, 6) (10, 12)
        8'b01000010, // Color (9, 8, 4) (11, 12)
        8'b00111110, // Color (12, 9, 6) (12, 12)
        8'b00111010, // Color (11, 9, 5) (13, 12)
        8'b00111110, // Color (12, 9, 6) (14, 12)
        8'b00111110, // Color (12, 9, 6) (15, 12)
        8'b00111100, // Color (10, 8, 5) (0, 13)
        8'b00111100, // Color (10, 8, 5) (1, 13)
        8'b00111010, // Color (11, 9, 5) (2, 13)
        8'b00111010, // Color (11, 9, 5) (3, 13)
        8'b01000010, // Color (9, 8, 4) (4, 13)
        8'b01000010, // Color (9, 8, 4) (5, 13)
        8'b00111100, // Color (10, 8, 5) (6, 13)
        8'b01000010, // Color (9, 8, 4) (7, 13)
        8'b01000010, // Color (9, 8, 4) (8, 13)
        8'b00111010, // Color (11, 9, 5) (9, 13)
        8'b00111010, // Color (11, 9, 5) (10, 13)
        8'b00111100, // Color (10, 8, 5) (11, 13)
        8'b00111010, // Color (11, 9, 5) (12, 13)
        8'b00111100, // Color (10, 8, 5) (13, 13)
        8'b00111100, // Color (10, 8, 5) (14, 13)
        8'b00111100, // Color (10, 8, 5) (15, 13)
        8'b00111100, // Color (10, 8, 5) (0, 14)
        8'b01000010, // Color (9, 8, 4) (1, 14)
        8'b01000010, // Color (9, 8, 4) (2, 14)
        8'b00111100, // Color (10, 8, 5) (3, 14)
        8'b00111010, // Color (11, 9, 5) (4, 14)
        8'b00111100, // Color (10, 8, 5) (5, 14)
        8'b01000010, // Color (9, 8, 4) (6, 14)
        8'b00110100, // Color (9, 7, 4) (7, 14)
        8'b00111010, // Color (11, 9, 5) (8, 14)
        8'b00111010, // Color (11, 9, 5) (9, 14)
        8'b00111100, // Color (10, 8, 5) (10, 14)
        8'b01000010, // Color (9, 8, 4) (11, 14)
        8'b01000010, // Color (9, 8, 4) (12, 14)
        8'b01000010, // Color (9, 8, 4) (13, 14)
        8'b01000010, // Color (9, 8, 4) (14, 14)
        8'b01000010, // Color (9, 8, 4) (15, 14)
        8'b01000100, // Color (6, 5, 2) (0, 15)
        8'b01000000, // Color (7, 6, 3) (1, 15)
        8'b01000000, // Color (7, 6, 3) (2, 15)
        8'b01000100, // Color (6, 5, 2) (3, 15)
        8'b01000100, // Color (6, 5, 2) (4, 15)
        8'b01000000, // Color (7, 6, 3) (5, 15)
        8'b00110100, // Color (9, 7, 4) (6, 15)
        8'b00110100, // Color (9, 7, 4) (7, 15)
        8'b00110100, // Color (9, 7, 4) (8, 15)
        8'b01000000, // Color (7, 6, 3) (9, 15)
        8'b01000100, // Color (6, 5, 2) (10, 15)
        8'b01000000, // Color (7, 6, 3) (11, 15)
        8'b01000100, // Color (6, 5, 2) (12, 15)
        8'b01000100, // Color (6, 5, 2) (13, 15)
        8'b01000100, // Color (6, 5, 2) (14, 15)
        8'b01000100, // Color (6, 5, 2) (15, 15)
        // 06_flowering_azalea_leaves
        8'b01000110, // Color (5, 6, 2) (0, 0)
        8'b01001000, // Color (0, 0, 0) (1, 0)
        8'b01001010, // Color (3, 4, 2) (2, 0)
        8'b01000110, // Color (5, 6, 2) (3, 0)
        8'b01000110, // Color (5, 6, 2) (4, 0)
        8'b01001100, // Color (6, 8, 3) (5, 0)
        8'b01001110, // Color (7, 9, 2) (6, 0)
        8'b01000110, // Color (5, 6, 2) (7, 0)
        8'b01000110, // Color (5, 6, 2) (8, 0)
        8'b01001000, // Color (0, 0, 0) (9, 0)
        8'b01001010, // Color (3, 4, 2) (10, 0)
        8'b01001010, // Color (3, 4, 2) (11, 0)
        8'b01001010, // Color (3, 4, 2) (12, 0)
        8'b01001000, // Color (0, 0, 0) (13, 0)
        8'b01000110, // Color (5, 6, 2) (14, 0)
        8'b01001100, // Color (6, 8, 3) (15, 0)
        8'b01001100, // Color (6, 8, 3) (0, 1)
        8'b01001000, // Color (0, 0, 0) (1, 1)
        8'b01001000, // Color (0, 0, 0) (2, 1)
        8'b01001010, // Color (3, 4, 2) (3, 1)
        8'b01001010, // Color (3, 4, 2) (4, 1)
        8'b01001110, // Color (7, 9, 2) (5, 1)
        8'b01001110, // Color (7, 9, 2) (6, 1)
        8'b01000110, // Color (5, 6, 2) (7, 1)
        8'b01000110, // Color (5, 6, 2) (8, 1)
        8'b01001000, // Color (0, 0, 0) (9, 1)
        8'b01001100, // Color (6, 8, 3) (10, 1)
        8'b01001100, // Color (6, 8, 3) (11, 1)
        8'b01001110, // Color (7, 9, 2) (12, 1)
        8'b01001000, // Color (0, 0, 0) (13, 1)
        8'b01001000, // Color (0, 0, 0) (14, 1)
        8'b01001100, // Color (6, 8, 3) (15, 1)
        8'b01001010, // Color (3, 4, 2) (0, 2)
        8'b01001000, // Color (0, 0, 0) (1, 2)
        8'b01000110, // Color (5, 6, 2) (2, 2)
        8'b01000110, // Color (5, 6, 2) (3, 2)
        8'b01000110, // Color (5, 6, 2) (4, 2)
        8'b01000110, // Color (5, 6, 2) (5, 2)
        8'b01001000, // Color (0, 0, 0) (6, 2)
        8'b01001000, // Color (0, 0, 0) (7, 2)
        8'b01001110, // Color (7, 9, 2) (8, 2)
        8'b01001100, // Color (6, 8, 3) (9, 2)
        8'b01001100, // Color (6, 8, 3) (10, 2)
        8'b01010000, // Color (11, 6, 12) (11, 2)
        8'b01010010, // Color (13, 7, 14) (12, 2)
        8'b01010000, // Color (11, 6, 12) (13, 2)
        8'b01001000, // Color (0, 0, 0) (14, 2)
        8'b01001010, // Color (3, 4, 2) (15, 2)
        8'b01001110, // Color (7, 9, 2) (0, 3)
        8'b01001100, // Color (6, 8, 3) (1, 3)
        8'b01000110, // Color (5, 6, 2) (2, 3)
        8'b01001110, // Color (7, 9, 2) (3, 3)
        8'b01001100, // Color (6, 8, 3) (4, 3)
        8'b01000110, // Color (5, 6, 2) (5, 3)
        8'b01001010, // Color (3, 4, 2) (6, 3)
        8'b01001000, // Color (0, 0, 0) (7, 3)
        8'b01001110, // Color (7, 9, 2) (8, 3)
        8'b01001110, // Color (7, 9, 2) (9, 3)
        8'b01000110, // Color (5, 6, 2) (10, 3)
        8'b01010010, // Color (13, 7, 14) (11, 3)
        8'b01001010, // Color (3, 4, 2) (12, 3)
        8'b01010010, // Color (13, 7, 14) (13, 3)
        8'b01001000, // Color (0, 0, 0) (14, 3)
        8'b01001010, // Color (3, 4, 2) (15, 3)
        8'b01001110, // Color (7, 9, 2) (0, 4)
        8'b01001110, // Color (7, 9, 2) (1, 4)
        8'b01001000, // Color (0, 0, 0) (2, 4)
        8'b01001110, // Color (7, 9, 2) (3, 4)
        8'b01001110, // Color (7, 9, 2) (4, 4)
        8'b01001010, // Color (3, 4, 2) (5, 4)
        8'b01001010, // Color (3, 4, 2) (6, 4)
        8'b01001000, // Color (0, 0, 0) (7, 4)
        8'b01001010, // Color (3, 4, 2) (8, 4)
        8'b01000110, // Color (5, 6, 2) (9, 4)
        8'b01000110, // Color (5, 6, 2) (10, 4)
        8'b01010000, // Color (11, 6, 12) (11, 4)
        8'b01010010, // Color (13, 7, 14) (12, 4)
        8'b01010100, // Color (9, 5, 8) (13, 4)
        8'b01001000, // Color (0, 0, 0) (14, 4)
        8'b01001000, // Color (0, 0, 0) (15, 4)
        8'b01001000, // Color (0, 0, 0) (0, 5)
        8'b01001000, // Color (0, 0, 0) (1, 5)
        8'b01001000, // Color (0, 0, 0) (2, 5)
        8'b01000110, // Color (5, 6, 2) (3, 5)
        8'b01000110, // Color (5, 6, 2) (4, 5)
        8'b01001010, // Color (3, 4, 2) (5, 5)
        8'b01001000, // Color (0, 0, 0) (6, 5)
        8'b01001010, // Color (3, 4, 2) (7, 5)
        8'b01001010, // Color (3, 4, 2) (8, 5)
        8'b01001010, // Color (3, 4, 2) (9, 5)
        8'b01001000, // Color (0, 0, 0) (10, 5)
        8'b01001000, // Color (0, 0, 0) (11, 5)
        8'b01001110, // Color (7, 9, 2) (12, 5)
        8'b01001110, // Color (7, 9, 2) (13, 5)
        8'b01001100, // Color (6, 8, 3) (14, 5)
        8'b01001100, // Color (6, 8, 3) (15, 5)
        8'b01001110, // Color (7, 9, 2) (0, 6)
        8'b01000110, // Color (5, 6, 2) (1, 6)
        8'b01001010, // Color (3, 4, 2) (2, 6)
        8'b01001000, // Color (0, 0, 0) (3, 6)
        8'b01001000, // Color (0, 0, 0) (4, 6)
        8'b01001000, // Color (0, 0, 0) (5, 6)
        8'b01001100, // Color (6, 8, 3) (6, 6)
        8'b01001110, // Color (7, 9, 2) (7, 6)
        8'b01001110, // Color (7, 9, 2) (8, 6)
        8'b01001110, // Color (7, 9, 2) (9, 6)
        8'b01000110, // Color (5, 6, 2) (10, 6)
        8'b01001010, // Color (3, 4, 2) (11, 6)
        8'b01001000, // Color (0, 0, 0) (12, 6)
        8'b01000110, // Color (5, 6, 2) (13, 6)
        8'b01001100, // Color (6, 8, 3) (14, 6)
        8'b01001100, // Color (6, 8, 3) (15, 6)
        8'b01001110, // Color (7, 9, 2) (0, 7)
        8'b01010000, // Color (11, 6, 12) (1, 7)
        8'b01010010, // Color (13, 7, 14) (2, 7)
        8'b01010100, // Color (9, 5, 8) (3, 7)
        8'b01001000, // Color (0, 0, 0) (4, 7)
        8'b01001000, // Color (0, 0, 0) (5, 7)
        8'b01000110, // Color (5, 6, 2) (6, 7)
        8'b01001110, // Color (7, 9, 2) (7, 7)
        8'b01001110, // Color (7, 9, 2) (8, 7)
        8'b01001110, // Color (7, 9, 2) (9, 7)
        8'b01001100, // Color (6, 8, 3) (10, 7)
        8'b01001010, // Color (3, 4, 2) (11, 7)
        8'b01001010, // Color (3, 4, 2) (12, 7)
        8'b01000110, // Color (5, 6, 2) (13, 7)
        8'b01000110, // Color (5, 6, 2) (14, 7)
        8'b01001110, // Color (7, 9, 2) (15, 7)
        8'b01001010, // Color (3, 4, 2) (0, 8)
        8'b01010010, // Color (13, 7, 14) (1, 8)
        8'b01001010, // Color (3, 4, 2) (2, 8)
        8'b01010000, // Color (11, 6, 12) (3, 8)
        8'b01001100, // Color (6, 8, 3) (4, 8)
        8'b01000110, // Color (5, 6, 2) (5, 8)
        8'b01001100, // Color (6, 8, 3) (6, 8)
        8'b01000110, // Color (5, 6, 2) (7, 8)
        8'b01000110, // Color (5, 6, 2) (8, 8)
        8'b01001110, // Color (7, 9, 2) (9, 8)
        8'b01001110, // Color (7, 9, 2) (10, 8)
        8'b01000110, // Color (5, 6, 2) (11, 8)
        8'b01001010, // Color (3, 4, 2) (12, 8)
        8'b01001010, // Color (3, 4, 2) (13, 8)
        8'b01000110, // Color (5, 6, 2) (14, 8)
        8'b01000110, // Color (5, 6, 2) (15, 8)
        8'b01000110, // Color (5, 6, 2) (0, 9)
        8'b01010100, // Color (9, 5, 8) (1, 9)
        8'b01010000, // Color (11, 6, 12) (2, 9)
        8'b01010100, // Color (9, 5, 8) (3, 9)
        8'b01001110, // Color (7, 9, 2) (4, 9)
        8'b01000110, // Color (5, 6, 2) (5, 9)
        8'b01001110, // Color (7, 9, 2) (6, 9)
        8'b01001100, // Color (6, 8, 3) (7, 9)
        8'b01000110, // Color (5, 6, 2) (8, 9)
        8'b01001110, // Color (7, 9, 2) (9, 9)
        8'b01001100, // Color (6, 8, 3) (10, 9)
        8'b01001100, // Color (6, 8, 3) (11, 9)
        8'b01001110, // Color (7, 9, 2) (12, 9)
        8'b01001000, // Color (0, 0, 0) (13, 9)
        8'b01001100, // Color (6, 8, 3) (14, 9)
        8'b01001100, // Color (6, 8, 3) (15, 9)
        8'b01001100, // Color (6, 8, 3) (0, 10)
        8'b01000110, // Color (5, 6, 2) (1, 10)
        8'b01000110, // Color (5, 6, 2) (2, 10)
        8'b01001110, // Color (7, 9, 2) (3, 10)
        8'b01000110, // Color (5, 6, 2) (4, 10)
        8'b01001000, // Color (0, 0, 0) (5, 10)
        8'b01001110, // Color (7, 9, 2) (6, 10)
        8'b01001110, // Color (7, 9, 2) (7, 10)
        8'b01001100, // Color (6, 8, 3) (8, 10)
        8'b01001000, // Color (0, 0, 0) (9, 10)
        8'b01001000, // Color (0, 0, 0) (10, 10)
        8'b01001110, // Color (7, 9, 2) (11, 10)
        8'b01001110, // Color (7, 9, 2) (12, 10)
        8'b01001000, // Color (0, 0, 0) (13, 10)
        8'b01001100, // Color (6, 8, 3) (14, 10)
        8'b01001100, // Color (6, 8, 3) (15, 10)
        8'b01001100, // Color (6, 8, 3) (0, 11)
        8'b01001000, // Color (0, 0, 0) (1, 11)
        8'b01001000, // Color (0, 0, 0) (2, 11)
        8'b01001010, // Color (3, 4, 2) (3, 11)
        8'b01001010, // Color (3, 4, 2) (4, 11)
        8'b01000110, // Color (5, 6, 2) (5, 11)
        8'b01001100, // Color (6, 8, 3) (6, 11)
        8'b01000110, // Color (5, 6, 2) (7, 11)
        8'b01001000, // Color (0, 0, 0) (8, 11)
        8'b01010100, // Color (9, 5, 8) (9, 11)
        8'b01010000, // Color (11, 6, 12) (10, 11)
        8'b01010100, // Color (9, 5, 8) (11, 11)
        8'b01000110, // Color (5, 6, 2) (12, 11)
        8'b01000110, // Color (5, 6, 2) (13, 11)
        8'b01001000, // Color (0, 0, 0) (14, 11)
        8'b01001100, // Color (6, 8, 3) (15, 11)
        8'b01001000, // Color (0, 0, 0) (0, 12)
        8'b01001010, // Color (3, 4, 2) (1, 12)
        8'b01000110, // Color (5, 6, 2) (2, 12)
        8'b01000110, // Color (5, 6, 2) (3, 12)
        8'b01001010, // Color (3, 4, 2) (4, 12)
        8'b01000110, // Color (5, 6, 2) (5, 12)
        8'b01000110, // Color (5, 6, 2) (6, 12)
        8'b01001000, // Color (0, 0, 0) (7, 12)
        8'b01000110, // Color (5, 6, 2) (8, 12)
        8'b01010000, // Color (11, 6, 12) (9, 12)
        8'b01001010, // Color (3, 4, 2) (10, 12)
        8'b01010000, // Color (11, 6, 12) (11, 12)
        8'b01001100, // Color (6, 8, 3) (12, 12)
        8'b01000110, // Color (5, 6, 2) (13, 12)
        8'b01001010, // Color (3, 4, 2) (14, 12)
        8'b01001010, // Color (3, 4, 2) (15, 12)
        8'b01001000, // Color (0, 0, 0) (0, 13)
        8'b01001100, // Color (6, 8, 3) (1, 13)
        8'b01001100, // Color (6, 8, 3) (2, 13)
        8'b01001110, // Color (7, 9, 2) (3, 13)
        8'b01001100, // Color (6, 8, 3) (4, 13)
        8'b01001100, // Color (6, 8, 3) (5, 13)
        8'b01001010, // Color (3, 4, 2) (6, 13)
        8'b01001000, // Color (0, 0, 0) (7, 13)
        8'b01000110, // Color (5, 6, 2) (8, 13)
        8'b01010100, // Color (9, 5, 8) (9, 13)
        8'b01010000, // Color (11, 6, 12) (10, 13)
        8'b01010100, // Color (9, 5, 8) (11, 13)
        8'b01001100, // Color (6, 8, 3) (12, 13)
        8'b01000110, // Color (5, 6, 2) (13, 13)
        8'b01001010, // Color (3, 4, 2) (14, 13)
        8'b01001010, // Color (3, 4, 2) (15, 13)
        8'b01000110, // Color (5, 6, 2) (0, 14)
        8'b01001100, // Color (6, 8, 3) (1, 14)
        8'b01001110, // Color (7, 9, 2) (2, 14)
        8'b01001100, // Color (6, 8, 3) (3, 14)
        8'b01001110, // Color (7, 9, 2) (4, 14)
        8'b01001100, // Color (6, 8, 3) (5, 14)
        8'b01001010, // Color (3, 4, 2) (6, 14)
        8'b01001010, // Color (3, 4, 2) (7, 14)
        8'b01001000, // Color (0, 0, 0) (8, 14)
        8'b01001000, // Color (0, 0, 0) (9, 14)
        8'b01000110, // Color (5, 6, 2) (10, 14)
        8'b01000110, // Color (5, 6, 2) (11, 14)
        8'b01001010, // Color (3, 4, 2) (12, 14)
        8'b01001100, // Color (6, 8, 3) (13, 14)
        8'b01001100, // Color (6, 8, 3) (14, 14)
        8'b01001000, // Color (0, 0, 0) (15, 14)
        8'b01000110, // Color (5, 6, 2) (0, 15)
        8'b01000110, // Color (5, 6, 2) (1, 15)
        8'b01000110, // Color (5, 6, 2) (2, 15)
        8'b01001110, // Color (7, 9, 2) (3, 15)
        8'b01001110, // Color (7, 9, 2) (4, 15)
        8'b01001000, // Color (0, 0, 0) (5, 15)
        8'b01001000, // Color (0, 0, 0) (6, 15)
        8'b01001010, // Color (3, 4, 2) (7, 15)
        8'b01001000, // Color (0, 0, 0) (8, 15)
        8'b01001000, // Color (0, 0, 0) (9, 15)
        8'b01001000, // Color (0, 0, 0) (10, 15)
        8'b01001010, // Color (3, 4, 2) (11, 15)
        8'b01001010, // Color (3, 4, 2) (12, 15)
        8'b01001100, // Color (6, 8, 3) (13, 15)
        8'b01001100, // Color (6, 8, 3) (14, 15)
        8'b01000110, // Color (5, 6, 2) (15, 15)
        // 07_jukebox_side
        8'b01010110, // Color (2, 2, 2) (0, 0)
        8'b01010110, // Color (2, 2, 2) (1, 0)
        8'b01010110, // Color (2, 2, 2) (2, 0)
        8'b01010110, // Color (2, 2, 2) (3, 0)
        8'b01010110, // Color (2, 2, 2) (4, 0)
        8'b01010110, // Color (2, 2, 2) (5, 0)
        8'b01010110, // Color (2, 2, 2) (6, 0)
        8'b01010110, // Color (2, 2, 2) (7, 0)
        8'b01010110, // Color (2, 2, 2) (8, 0)
        8'b01010110, // Color (2, 2, 2) (9, 0)
        8'b01010110, // Color (2, 2, 2) (10, 0)
        8'b01010110, // Color (2, 2, 2) (11, 0)
        8'b01010110, // Color (2, 2, 2) (12, 0)
        8'b01010110, // Color (2, 2, 2) (13, 0)
        8'b01010110, // Color (2, 2, 2) (14, 0)
        8'b01010110, // Color (2, 2, 2) (15, 0)
        8'b01010110, // Color (2, 2, 2) (0, 1)
        8'b00001000, // Color (5, 3, 2) (1, 1)
        8'b00000110, // Color (7, 5, 3) (2, 1)
        8'b01011000, // Color (9, 5, 4) (3, 1)
        8'b01011000, // Color (9, 5, 4) (4, 1)
        8'b00000110, // Color (7, 5, 3) (5, 1)
        8'b00000110, // Color (7, 5, 3) (6, 1)
        8'b01011000, // Color (9, 5, 4) (7, 1)
        8'b01011000, // Color (9, 5, 4) (8, 1)
        8'b01011000, // Color (9, 5, 4) (9, 1)
        8'b01011000, // Color (9, 5, 4) (10, 1)
        8'b00000110, // Color (7, 5, 3) (11, 1)
        8'b01011000, // Color (9, 5, 4) (12, 1)
        8'b00000110, // Color (7, 5, 3) (13, 1)
        8'b00001000, // Color (5, 3, 2) (14, 1)
        8'b01010110, // Color (2, 2, 2) (15, 1)
        8'b01010110, // Color (2, 2, 2) (0, 2)
        8'b00000110, // Color (7, 5, 3) (1, 2)
        8'b01011000, // Color (9, 5, 4) (2, 2)
        8'b01011010, // Color (4, 2, 1) (3, 2)
        8'b01011000, // Color (9, 5, 4) (4, 2)
        8'b01011010, // Color (4, 2, 1) (5, 2)
        8'b01011000, // Color (9, 5, 4) (6, 2)
        8'b01011010, // Color (4, 2, 1) (7, 2)
        8'b01011000, // Color (9, 5, 4) (8, 2)
        8'b01011010, // Color (4, 2, 1) (9, 2)
        8'b01011000, // Color (9, 5, 4) (10, 2)
        8'b01011010, // Color (4, 2, 1) (11, 2)
        8'b00000110, // Color (7, 5, 3) (12, 2)
        8'b01011010, // Color (4, 2, 1) (13, 2)
        8'b00000110, // Color (7, 5, 3) (14, 2)
        8'b01010110, // Color (2, 2, 2) (15, 2)
        8'b01010110, // Color (2, 2, 2) (0, 3)
        8'b01011000, // Color (9, 5, 4) (1, 3)
        8'b01011010, // Color (4, 2, 1) (2, 3)
        8'b01011000, // Color (9, 5, 4) (3, 3)
        8'b00001000, // Color (5, 3, 2) (4, 3)
        8'b01011010, // Color (4, 2, 1) (5, 3)
        8'b00001000, // Color (5, 3, 2) (6, 3)
        8'b01011000, // Color (9, 5, 4) (7, 3)
        8'b00001000, // Color (5, 3, 2) (8, 3)
        8'b01011010, // Color (4, 2, 1) (9, 3)
        8'b00001000, // Color (5, 3, 2) (10, 3)
        8'b01011000, // Color (9, 5, 4) (11, 3)
        8'b00001000, // Color (5, 3, 2) (12, 3)
        8'b01011010, // Color (4, 2, 1) (13, 3)
        8'b01011000, // Color (9, 5, 4) (14, 3)
        8'b01010110, // Color (2, 2, 2) (15, 3)
        8'b01010110, // Color (2, 2, 2) (0, 4)
        8'b01011000, // Color (9, 5, 4) (1, 4)
        8'b01011000, // Color (9, 5, 4) (2, 4)
        8'b01011010, // Color (4, 2, 1) (3, 4)
        8'b01011000, // Color (9, 5, 4) (4, 4)
        8'b00001000, // Color (5, 3, 2) (5, 4)
        8'b01011000, // Color (9, 5, 4) (6, 4)
        8'b01011010, // Color (4, 2, 1) (7, 4)
        8'b01011000, // Color (9, 5, 4) (8, 4)
        8'b00001000, // Color (5, 3, 2) (9, 4)
        8'b01011000, // Color (9, 5, 4) (10, 4)
        8'b01011010, // Color (4, 2, 1) (11, 4)
        8'b00000110, // Color (7, 5, 3) (12, 4)
        8'b00001000, // Color (5, 3, 2) (13, 4)
        8'b01011000, // Color (9, 5, 4) (14, 4)
        8'b01010110, // Color (2, 2, 2) (15, 4)
        8'b01010110, // Color (2, 2, 2) (0, 5)
        8'b00000110, // Color (7, 5, 3) (1, 5)
        8'b00001000, // Color (5, 3, 2) (2, 5)
        8'b01011010, // Color (4, 2, 1) (3, 5)
        8'b00001000, // Color (5, 3, 2) (4, 5)
        8'b01011000, // Color (9, 5, 4) (5, 5)
        8'b00001000, // Color (5, 3, 2) (6, 5)
        8'b01011010, // Color (4, 2, 1) (7, 5)
        8'b00001000, // Color (5, 3, 2) (8, 5)
        8'b01011000, // Color (9, 5, 4) (9, 5)
        8'b00001000, // Color (5, 3, 2) (10, 5)
        8'b01011010, // Color (4, 2, 1) (11, 5)
        8'b00001000, // Color (5, 3, 2) (12, 5)
        8'b00000110, // Color (7, 5, 3) (13, 5)
        8'b01011000, // Color (9, 5, 4) (14, 5)
        8'b01010110, // Color (2, 2, 2) (15, 5)
        8'b01010110, // Color (2, 2, 2) (0, 6)
        8'b01011000, // Color (9, 5, 4) (1, 6)
        8'b01011000, // Color (9, 5, 4) (2, 6)
        8'b00001000, // Color (5, 3, 2) (3, 6)
        8'b01011000, // Color (9, 5, 4) (4, 6)
        8'b01011010, // Color (4, 2, 1) (5, 6)
        8'b01011000, // Color (9, 5, 4) (6, 6)
        8'b00001000, // Color (5, 3, 2) (7, 6)
        8'b00000110, // Color (7, 5, 3) (8, 6)
        8'b01011010, // Color (4, 2, 1) (9, 6)
        8'b01011000, // Color (9, 5, 4) (10, 6)
        8'b00001000, // Color (5, 3, 2) (11, 6)
        8'b00000110, // Color (7, 5, 3) (12, 6)
        8'b01011010, // Color (4, 2, 1) (13, 6)
        8'b00000110, // Color (7, 5, 3) (14, 6)
        8'b01010110, // Color (2, 2, 2) (15, 6)
        8'b01010110, // Color (2, 2, 2) (0, 7)
        8'b00000110, // Color (7, 5, 3) (1, 7)
        8'b01011010, // Color (4, 2, 1) (2, 7)
        8'b01011000, // Color (9, 5, 4) (3, 7)
        8'b00001000, // Color (5, 3, 2) (4, 7)
        8'b01011010, // Color (4, 2, 1) (5, 7)
        8'b00001000, // Color (5, 3, 2) (6, 7)
        8'b01011000, // Color (9, 5, 4) (7, 7)
        8'b00001000, // Color (5, 3, 2) (8, 7)
        8'b01011010, // Color (4, 2, 1) (9, 7)
        8'b00001000, // Color (5, 3, 2) (10, 7)
        8'b01011000, // Color (9, 5, 4) (11, 7)
        8'b00001000, // Color (5, 3, 2) (12, 7)
        8'b01011010, // Color (4, 2, 1) (13, 7)
        8'b00001000, // Color (5, 3, 2) (14, 7)
        8'b01010110, // Color (2, 2, 2) (15, 7)
        8'b01010110, // Color (2, 2, 2) (0, 8)
        8'b00001000, // Color (5, 3, 2) (1, 8)
        8'b00000110, // Color (7, 5, 3) (2, 8)
        8'b01011010, // Color (4, 2, 1) (3, 8)
        8'b01011000, // Color (9, 5, 4) (4, 8)
        8'b00001000, // Color (5, 3, 2) (5, 8)
        8'b00000110, // Color (7, 5, 3) (6, 8)
        8'b01011010, // Color (4, 2, 1) (7, 8)
        8'b01011000, // Color (9, 5, 4) (8, 8)
        8'b00001000, // Color (5, 3, 2) (9, 8)
        8'b00000110, // Color (7, 5, 3) (10, 8)
        8'b01011010, // Color (4, 2, 1) (11, 8)
        8'b00000110, // Color (7, 5, 3) (12, 8)
        8'b00001000, // Color (5, 3, 2) (13, 8)
        8'b01011000, // Color (9, 5, 4) (14, 8)
        8'b01010110, // Color (2, 2, 2) (15, 8)
        8'b01010110, // Color (2, 2, 2) (0, 9)
        8'b00000110, // Color (7, 5, 3) (1, 9)
        8'b00001000, // Color (5, 3, 2) (2, 9)
        8'b01011010, // Color (4, 2, 1) (3, 9)
        8'b00001000, // Color (5, 3, 2) (4, 9)
        8'b01011000, // Color (9, 5, 4) (5, 9)
        8'b00001000, // Color (5, 3, 2) (6, 9)
        8'b01011010, // Color (4, 2, 1) (7, 9)
        8'b00001000, // Color (5, 3, 2) (8, 9)
        8'b01011000, // Color (9, 5, 4) (9, 9)
        8'b00001000, // Color (5, 3, 2) (10, 9)
        8'b01011010, // Color (4, 2, 1) (11, 9)
        8'b00001000, // Color (5, 3, 2) (12, 9)
        8'b00000110, // Color (7, 5, 3) (13, 9)
        8'b00000110, // Color (7, 5, 3) (14, 9)
        8'b01010110, // Color (2, 2, 2) (15, 9)
        8'b01010110, // Color (2, 2, 2) (0, 10)
        8'b01011000, // Color (9, 5, 4) (1, 10)
        8'b00000110, // Color (7, 5, 3) (2, 10)
        8'b00001000, // Color (5, 3, 2) (3, 10)
        8'b00000110, // Color (7, 5, 3) (4, 10)
        8'b01011010, // Color (4, 2, 1) (5, 10)
        8'b01011000, // Color (9, 5, 4) (6, 10)
        8'b00001000, // Color (5, 3, 2) (7, 10)
        8'b00000110, // Color (7, 5, 3) (8, 10)
        8'b01011010, // Color (4, 2, 1) (9, 10)
        8'b01011000, // Color (9, 5, 4) (10, 10)
        8'b00001000, // Color (5, 3, 2) (11, 10)
        8'b00000110, // Color (7, 5, 3) (12, 10)
        8'b01011010, // Color (4, 2, 1) (13, 10)
        8'b00000110, // Color (7, 5, 3) (14, 10)
        8'b01010110, // Color (2, 2, 2) (15, 10)
        8'b01010110, // Color (2, 2, 2) (0, 11)
        8'b00000110, // Color (7, 5, 3) (1, 11)
        8'b01011010, // Color (4, 2, 1) (2, 11)
        8'b00000110, // Color (7, 5, 3) (3, 11)
        8'b00001000, // Color (5, 3, 2) (4, 11)
        8'b01011010, // Color (4, 2, 1) (5, 11)
        8'b00001000, // Color (5, 3, 2) (6, 11)
        8'b00000110, // Color (7, 5, 3) (7, 11)
        8'b00001000, // Color (5, 3, 2) (8, 11)
        8'b01011010, // Color (4, 2, 1) (9, 11)
        8'b00001000, // Color (5, 3, 2) (10, 11)
        8'b00000110, // Color (7, 5, 3) (11, 11)
        8'b00001000, // Color (5, 3, 2) (12, 11)
        8'b01011010, // Color (4, 2, 1) (13, 11)
        8'b00001000, // Color (5, 3, 2) (14, 11)
        8'b01010110, // Color (2, 2, 2) (15, 11)
        8'b01010110, // Color (2, 2, 2) (0, 12)
        8'b00000110, // Color (7, 5, 3) (1, 12)
        8'b00001000, // Color (5, 3, 2) (2, 12)
        8'b01011010, // Color (4, 2, 1) (3, 12)
        8'b00000110, // Color (7, 5, 3) (4, 12)
        8'b00001000, // Color (5, 3, 2) (5, 12)
        8'b00000110, // Color (7, 5, 3) (6, 12)
        8'b01011010, // Color (4, 2, 1) (7, 12)
        8'b00000110, // Color (7, 5, 3) (8, 12)
        8'b00001000, // Color (5, 3, 2) (9, 12)
        8'b00000110, // Color (7, 5, 3) (10, 12)
        8'b01011010, // Color (4, 2, 1) (11, 12)
        8'b00000110, // Color (7, 5, 3) (12, 12)
        8'b01011010, // Color (4, 2, 1) (13, 12)
        8'b00000110, // Color (7, 5, 3) (14, 12)
        8'b01010110, // Color (2, 2, 2) (15, 12)
        8'b01010110, // Color (2, 2, 2) (0, 13)
        8'b00001000, // Color (5, 3, 2) (1, 13)
        8'b01011010, // Color (4, 2, 1) (2, 13)
        8'b01011010, // Color (4, 2, 1) (3, 13)
        8'b01011010, // Color (4, 2, 1) (4, 13)
        8'b00000110, // Color (7, 5, 3) (5, 13)
        8'b01011010, // Color (4, 2, 1) (6, 13)
        8'b01011010, // Color (4, 2, 1) (7, 13)
        8'b01011010, // Color (4, 2, 1) (8, 13)
        8'b00000110, // Color (7, 5, 3) (9, 13)
        8'b01011010, // Color (4, 2, 1) (10, 13)
        8'b01011010, // Color (4, 2, 1) (11, 13)
        8'b01011010, // Color (4, 2, 1) (12, 13)
        8'b00000110, // Color (7, 5, 3) (13, 13)
        8'b00001000, // Color (5, 3, 2) (14, 13)
        8'b01010110, // Color (2, 2, 2) (15, 13)
        8'b01010110, // Color (2, 2, 2) (0, 14)
        8'b00001000, // Color (5, 3, 2) (1, 14)
        8'b00001000, // Color (5, 3, 2) (2, 14)
        8'b00001000, // Color (5, 3, 2) (3, 14)
        8'b00001000, // Color (5, 3, 2) (4, 14)
        8'b00001000, // Color (5, 3, 2) (5, 14)
        8'b00001000, // Color (5, 3, 2) (6, 14)
        8'b00001000, // Color (5, 3, 2) (7, 14)
        8'b00001000, // Color (5, 3, 2) (8, 14)
        8'b00001000, // Color (5, 3, 2) (9, 14)
        8'b00001000, // Color (5, 3, 2) (10, 14)
        8'b00001000, // Color (5, 3, 2) (11, 14)
        8'b00001000, // Color (5, 3, 2) (12, 14)
        8'b00001000, // Color (5, 3, 2) (13, 14)
        8'b00001000, // Color (5, 3, 2) (14, 14)
        8'b01010110, // Color (2, 2, 2) (15, 14)
        8'b01010110, // Color (2, 2, 2) (0, 15)
        8'b01010110, // Color (2, 2, 2) (1, 15)
        8'b01010110, // Color (2, 2, 2) (2, 15)
        8'b01010110, // Color (2, 2, 2) (3, 15)
        8'b01010110, // Color (2, 2, 2) (4, 15)
        8'b01010110, // Color (2, 2, 2) (5, 15)
        8'b01010110, // Color (2, 2, 2) (6, 15)
        8'b01010110, // Color (2, 2, 2) (7, 15)
        8'b01010110, // Color (2, 2, 2) (8, 15)
        8'b01010110, // Color (2, 2, 2) (9, 15)
        8'b01010110, // Color (2, 2, 2) (10, 15)
        8'b01010110, // Color (2, 2, 2) (11, 15)
        8'b01010110, // Color (2, 2, 2) (12, 15)
        8'b01010110, // Color (2, 2, 2) (13, 15)
        8'b01010110, // Color (2, 2, 2) (14, 15)
        8'b01010110, // Color (2, 2, 2) (15, 15)
        // 08_
        8'b00001010, // Color (8, 8, 8) (0, 0)
        8'b00001010, // Color (8, 8, 8) (1, 0)
        8'b00001010, // Color (8, 8, 8) (2, 0)
        8'b00001010, // Color (8, 8, 8) (3, 0)
        8'b01011100, // Color (7, 7, 7) (4, 0)
        8'b01011100, // Color (7, 7, 7) (5, 0)
        8'b01011100, // Color (7, 7, 7) (6, 0)
        8'b01011100, // Color (7, 7, 7) (7, 0)
        8'b01011100, // Color (7, 7, 7) (8, 0)
        8'b00001100, // Color (6, 6, 6) (9, 0)
        8'b01011100, // Color (7, 7, 7) (10, 0)
        8'b01011100, // Color (7, 7, 7) (11, 0)
        8'b01011100, // Color (7, 7, 7) (12, 0)
        8'b01011100, // Color (7, 7, 7) (13, 0)
        8'b01011100, // Color (7, 7, 7) (14, 0)
        8'b01011100, // Color (7, 7, 7) (15, 0)
        8'b01011100, // Color (7, 7, 7) (0, 1)
        8'b01011100, // Color (7, 7, 7) (1, 1)
        8'b01011100, // Color (7, 7, 7) (2, 1)
        8'b01011100, // Color (7, 7, 7) (3, 1)
        8'b01011100, // Color (7, 7, 7) (4, 1)
        8'b01011100, // Color (7, 7, 7) (5, 1)
        8'b01011100, // Color (7, 7, 7) (6, 1)
        8'b01011100, // Color (7, 7, 7) (7, 1)
        8'b01011100, // Color (7, 7, 7) (8, 1)
        8'b01011100, // Color (7, 7, 7) (9, 1)
        8'b01011100, // Color (7, 7, 7) (10, 1)
        8'b00001100, // Color (6, 6, 6) (11, 1)
        8'b00001100, // Color (6, 6, 6) (12, 1)
        8'b01011100, // Color (7, 7, 7) (13, 1)
        8'b01011100, // Color (7, 7, 7) (14, 1)
        8'b01011100, // Color (7, 7, 7) (15, 1)
        8'b01011100, // Color (7, 7, 7) (0, 2)
        8'b01011100, // Color (7, 7, 7) (1, 2)
        8'b00001100, // Color (6, 6, 6) (2, 2)
        8'b00001100, // Color (6, 6, 6) (3, 2)
        8'b01011100, // Color (7, 7, 7) (4, 2)
        8'b01011100, // Color (7, 7, 7) (5, 2)
        8'b01011100, // Color (7, 7, 7) (6, 2)
        8'b00001100, // Color (6, 6, 6) (7, 2)
        8'b01011100, // Color (7, 7, 7) (8, 2)
        8'b01011100, // Color (7, 7, 7) (9, 2)
        8'b01011100, // Color (7, 7, 7) (10, 2)
        8'b01011100, // Color (7, 7, 7) (11, 2)
        8'b01011100, // Color (7, 7, 7) (12, 2)
        8'b01011100, // Color (7, 7, 7) (13, 2)
        8'b01011100, // Color (7, 7, 7) (14, 2)
        8'b01011100, // Color (7, 7, 7) (15, 2)
        8'b01011100, // Color (7, 7, 7) (0, 3)
        8'b01011100, // Color (7, 7, 7) (1, 3)
        8'b00001010, // Color (8, 8, 8) (2, 3)
        8'b00001010, // Color (8, 8, 8) (3, 3)
        8'b01011100, // Color (7, 7, 7) (4, 3)
        8'b00001010, // Color (8, 8, 8) (5, 3)
        8'b01011100, // Color (7, 7, 7) (6, 3)
        8'b01011100, // Color (7, 7, 7) (7, 3)
        8'b00001010, // Color (8, 8, 8) (8, 3)
        8'b00001010, // Color (8, 8, 8) (9, 3)
        8'b01011100, // Color (7, 7, 7) (10, 3)
        8'b01011100, // Color (7, 7, 7) (11, 3)
        8'b01011100, // Color (7, 7, 7) (12, 3)
        8'b01011100, // Color (7, 7, 7) (13, 3)
        8'b01011100, // Color (7, 7, 7) (14, 3)
        8'b01011100, // Color (7, 7, 7) (15, 3)
        8'b01011100, // Color (7, 7, 7) (0, 4)
        8'b01011100, // Color (7, 7, 7) (1, 4)
        8'b01011100, // Color (7, 7, 7) (2, 4)
        8'b01011100, // Color (7, 7, 7) (3, 4)
        8'b01011100, // Color (7, 7, 7) (4, 4)
        8'b01011100, // Color (7, 7, 7) (5, 4)
        8'b01011100, // Color (7, 7, 7) (6, 4)
        8'b01011100, // Color (7, 7, 7) (7, 4)
        8'b01011100, // Color (7, 7, 7) (8, 4)
        8'b00001010, // Color (8, 8, 8) (9, 4)
        8'b00001010, // Color (8, 8, 8) (10, 4)
        8'b00001010, // Color (8, 8, 8) (11, 4)
        8'b00001010, // Color (8, 8, 8) (12, 4)
        8'b01011100, // Color (7, 7, 7) (13, 4)
        8'b01011100, // Color (7, 7, 7) (14, 4)
        8'b01011100, // Color (7, 7, 7) (15, 4)
        8'b01011100, // Color (7, 7, 7) (0, 5)
        8'b00001010, // Color (8, 8, 8) (1, 5)
        8'b01011100, // Color (7, 7, 7) (2, 5)
        8'b01011100, // Color (7, 7, 7) (3, 5)
        8'b01011100, // Color (7, 7, 7) (4, 5)
        8'b01011100, // Color (7, 7, 7) (5, 5)
        8'b01011100, // Color (7, 7, 7) (6, 5)
        8'b01011100, // Color (7, 7, 7) (7, 5)
        8'b01011100, // Color (7, 7, 7) (8, 5)
        8'b01011100, // Color (7, 7, 7) (9, 5)
        8'b01011100, // Color (7, 7, 7) (10, 5)
        8'b00001100, // Color (6, 6, 6) (11, 5)
        8'b01011100, // Color (7, 7, 7) (12, 5)
        8'b00001100, // Color (6, 6, 6) (13, 5)
        8'b01011100, // Color (7, 7, 7) (14, 5)
        8'b00001010, // Color (8, 8, 8) (15, 5)
        8'b01011100, // Color (7, 7, 7) (0, 6)
        8'b01011100, // Color (7, 7, 7) (1, 6)
        8'b01011100, // Color (7, 7, 7) (2, 6)
        8'b00001010, // Color (8, 8, 8) (3, 6)
        8'b00001010, // Color (8, 8, 8) (4, 6)
        8'b00001010, // Color (8, 8, 8) (5, 6)
        8'b01011100, // Color (7, 7, 7) (6, 6)
        8'b00001010, // Color (8, 8, 8) (7, 6)
        8'b00001010, // Color (8, 8, 8) (8, 6)
        8'b01011100, // Color (7, 7, 7) (9, 6)
        8'b01011100, // Color (7, 7, 7) (10, 6)
        8'b01011100, // Color (7, 7, 7) (11, 6)
        8'b01011100, // Color (7, 7, 7) (12, 6)
        8'b01011100, // Color (7, 7, 7) (13, 6)
        8'b01011100, // Color (7, 7, 7) (14, 6)
        8'b01011100, // Color (7, 7, 7) (15, 6)
        8'b01011100, // Color (7, 7, 7) (0, 7)
        8'b01011100, // Color (7, 7, 7) (1, 7)
        8'b00001100, // Color (6, 6, 6) (2, 7)
        8'b00001100, // Color (6, 6, 6) (3, 7)
        8'b01011100, // Color (7, 7, 7) (4, 7)
        8'b00001100, // Color (6, 6, 6) (5, 7)
        8'b01011100, // Color (7, 7, 7) (6, 7)
        8'b01011100, // Color (7, 7, 7) (7, 7)
        8'b01011100, // Color (7, 7, 7) (8, 7)
        8'b01011100, // Color (7, 7, 7) (9, 7)
        8'b01011100, // Color (7, 7, 7) (10, 7)
        8'b01011100, // Color (7, 7, 7) (11, 7)
        8'b01011100, // Color (7, 7, 7) (12, 7)
        8'b01011100, // Color (7, 7, 7) (13, 7)
        8'b01011100, // Color (7, 7, 7) (14, 7)
        8'b01011100, // Color (7, 7, 7) (15, 7)
        8'b00001010, // Color (8, 8, 8) (0, 8)
        8'b00001010, // Color (8, 8, 8) (1, 8)
        8'b00001010, // Color (8, 8, 8) (2, 8)
        8'b01011100, // Color (7, 7, 7) (3, 8)
        8'b00001010, // Color (8, 8, 8) (4, 8)
        8'b01011100, // Color (7, 7, 7) (5, 8)
        8'b01011100, // Color (7, 7, 7) (6, 8)
        8'b00001010, // Color (8, 8, 8) (7, 8)
        8'b00001010, // Color (8, 8, 8) (8, 8)
        8'b00001010, // Color (8, 8, 8) (9, 8)
        8'b01011100, // Color (7, 7, 7) (10, 8)
        8'b01011100, // Color (7, 7, 7) (11, 8)
        8'b01011100, // Color (7, 7, 7) (12, 8)
        8'b01011100, // Color (7, 7, 7) (13, 8)
        8'b01011100, // Color (7, 7, 7) (14, 8)
        8'b01011100, // Color (7, 7, 7) (15, 8)
        8'b01011100, // Color (7, 7, 7) (0, 9)
        8'b01011100, // Color (7, 7, 7) (1, 9)
        8'b00001010, // Color (8, 8, 8) (2, 9)
        8'b01011100, // Color (7, 7, 7) (3, 9)
        8'b01011100, // Color (7, 7, 7) (4, 9)
        8'b01011100, // Color (7, 7, 7) (5, 9)
        8'b00001010, // Color (8, 8, 8) (6, 9)
        8'b00001010, // Color (8, 8, 8) (7, 9)
        8'b00001010, // Color (8, 8, 8) (8, 9)
        8'b01011100, // Color (7, 7, 7) (9, 9)
        8'b01011100, // Color (7, 7, 7) (10, 9)
        8'b00001010, // Color (8, 8, 8) (11, 9)
        8'b00001010, // Color (8, 8, 8) (12, 9)
        8'b00001010, // Color (8, 8, 8) (13, 9)
        8'b00001010, // Color (8, 8, 8) (14, 9)
        8'b01011100, // Color (7, 7, 7) (15, 9)
        8'b00001100, // Color (6, 6, 6) (0, 10)
        8'b01011100, // Color (7, 7, 7) (1, 10)
        8'b01011100, // Color (7, 7, 7) (2, 10)
        8'b01011100, // Color (7, 7, 7) (3, 10)
        8'b01011100, // Color (7, 7, 7) (4, 10)
        8'b01011100, // Color (7, 7, 7) (5, 10)
        8'b00001100, // Color (6, 6, 6) (6, 10)
        8'b00001100, // Color (6, 6, 6) (7, 10)
        8'b01011100, // Color (7, 7, 7) (8, 10)
        8'b01011100, // Color (7, 7, 7) (9, 10)
        8'b01011100, // Color (7, 7, 7) (10, 10)
        8'b01011100, // Color (7, 7, 7) (11, 10)
        8'b01011100, // Color (7, 7, 7) (12, 10)
        8'b01011100, // Color (7, 7, 7) (13, 10)
        8'b01011100, // Color (7, 7, 7) (14, 10)
        8'b01011100, // Color (7, 7, 7) (15, 10)
        8'b01011100, // Color (7, 7, 7) (0, 11)
        8'b01011100, // Color (7, 7, 7) (1, 11)
        8'b01011100, // Color (7, 7, 7) (2, 11)
        8'b01011100, // Color (7, 7, 7) (3, 11)
        8'b01011100, // Color (7, 7, 7) (4, 11)
        8'b00001010, // Color (8, 8, 8) (5, 11)
        8'b00001010, // Color (8, 8, 8) (6, 11)
        8'b01011100, // Color (7, 7, 7) (7, 11)
        8'b01011100, // Color (7, 7, 7) (8, 11)
        8'b01011100, // Color (7, 7, 7) (9, 11)
        8'b01011100, // Color (7, 7, 7) (10, 11)
        8'b01011100, // Color (7, 7, 7) (11, 11)
        8'b00001010, // Color (8, 8, 8) (12, 11)
        8'b00001010, // Color (8, 8, 8) (13, 11)
        8'b01011100, // Color (7, 7, 7) (14, 11)
        8'b00001010, // Color (8, 8, 8) (15, 11)
        8'b01011100, // Color (7, 7, 7) (0, 12)
        8'b01011100, // Color (7, 7, 7) (1, 12)
        8'b01011100, // Color (7, 7, 7) (2, 12)
        8'b01011100, // Color (7, 7, 7) (3, 12)
        8'b01011100, // Color (7, 7, 7) (4, 12)
        8'b00001010, // Color (8, 8, 8) (5, 12)
        8'b01011100, // Color (7, 7, 7) (6, 12)
        8'b01011100, // Color (7, 7, 7) (7, 12)
        8'b01011100, // Color (7, 7, 7) (8, 12)
        8'b01011100, // Color (7, 7, 7) (9, 12)
        8'b01011100, // Color (7, 7, 7) (10, 12)
        8'b00001100, // Color (6, 6, 6) (11, 12)
        8'b00001100, // Color (6, 6, 6) (12, 12)
        8'b01011100, // Color (7, 7, 7) (13, 12)
        8'b00001100, // Color (6, 6, 6) (14, 12)
        8'b01011100, // Color (7, 7, 7) (15, 12)
        8'b00001010, // Color (8, 8, 8) (0, 13)
        8'b00001010, // Color (8, 8, 8) (1, 13)
        8'b01011100, // Color (7, 7, 7) (2, 13)
        8'b01011100, // Color (7, 7, 7) (3, 13)
        8'b01011100, // Color (7, 7, 7) (4, 13)
        8'b01011100, // Color (7, 7, 7) (5, 13)
        8'b01011100, // Color (7, 7, 7) (6, 13)
        8'b01011100, // Color (7, 7, 7) (7, 13)
        8'b01011100, // Color (7, 7, 7) (8, 13)
        8'b01011100, // Color (7, 7, 7) (9, 13)
        8'b01011100, // Color (7, 7, 7) (10, 13)
        8'b01011100, // Color (7, 7, 7) (11, 13)
        8'b01011100, // Color (7, 7, 7) (12, 13)
        8'b01011100, // Color (7, 7, 7) (13, 13)
        8'b01011100, // Color (7, 7, 7) (14, 13)
        8'b00001010, // Color (8, 8, 8) (15, 13)
        8'b01011100, // Color (7, 7, 7) (0, 14)
        8'b01011100, // Color (7, 7, 7) (1, 14)
        8'b01011100, // Color (7, 7, 7) (2, 14)
        8'b01011100, // Color (7, 7, 7) (3, 14)
        8'b01011100, // Color (7, 7, 7) (4, 14)
        8'b01011100, // Color (7, 7, 7) (5, 14)
        8'b01011100, // Color (7, 7, 7) (6, 14)
        8'b01011100, // Color (7, 7, 7) (7, 14)
        8'b01011100, // Color (7, 7, 7) (8, 14)
        8'b01011100, // Color (7, 7, 7) (9, 14)
        8'b01011100, // Color (7, 7, 7) (10, 14)
        8'b01011100, // Color (7, 7, 7) (11, 14)
        8'b00001010, // Color (8, 8, 8) (12, 14)
        8'b00001010, // Color (8, 8, 8) (13, 14)
        8'b00001010, // Color (8, 8, 8) (14, 14)
        8'b00001010, // Color (8, 8, 8) (15, 14)
        8'b01011100, // Color (7, 7, 7) (0, 15)
        8'b01011100, // Color (7, 7, 7) (1, 15)
        8'b01011100, // Color (7, 7, 7) (2, 15)
        8'b01011100, // Color (7, 7, 7) (3, 15)
        8'b01011100, // Color (7, 7, 7) (4, 15)
        8'b01011100, // Color (7, 7, 7) (5, 15)
        8'b01011100, // Color (7, 7, 7) (6, 15)
        8'b01011100, // Color (7, 7, 7) (7, 15)
        8'b01011100, // Color (7, 7, 7) (8, 15)
        8'b00001010, // Color (8, 8, 8) (9, 15)
        8'b00001010, // Color (8, 8, 8) (10, 15)
        8'b01011100, // Color (7, 7, 7) (11, 15)
        8'b01011100, // Color (7, 7, 7) (12, 15)
        8'b01011100, // Color (7, 7, 7) (13, 15)
        8'b01011100, // Color (7, 7, 7) (14, 15)
        8'b01011100, // Color (7, 7, 7) (15, 15)
        // 09_jukebox_top
        8'b01010110, // Color (2, 2, 2) (0, 0)
        8'b01010110, // Color (2, 2, 2) (1, 0)
        8'b01011110, // Color (3, 2, 2) (2, 0)
        8'b01011110, // Color (3, 2, 2) (3, 0)
        8'b01010110, // Color (2, 2, 2) (4, 0)
        8'b01010110, // Color (2, 2, 2) (5, 0)
        8'b01011110, // Color (3, 2, 2) (6, 0)
        8'b01011110, // Color (3, 2, 2) (7, 0)
        8'b01011110, // Color (3, 2, 2) (8, 0)
        8'b01011110, // Color (3, 2, 2) (9, 0)
        8'b01011110, // Color (3, 2, 2) (10, 0)
        8'b01010110, // Color (2, 2, 2) (11, 0)
        8'b01011110, // Color (3, 2, 2) (12, 0)
        8'b01010110, // Color (2, 2, 2) (13, 0)
        8'b01010110, // Color (2, 2, 2) (14, 0)
        8'b01010110, // Color (2, 2, 2) (15, 0)
        8'b01010110, // Color (2, 2, 2) (0, 1)
        8'b00001000, // Color (5, 3, 2) (1, 1)
        8'b00001000, // Color (5, 3, 2) (2, 1)
        8'b00000110, // Color (7, 5, 3) (3, 1)
        8'b00000110, // Color (7, 5, 3) (4, 1)
        8'b00001000, // Color (5, 3, 2) (5, 1)
        8'b00001000, // Color (5, 3, 2) (6, 1)
        8'b00001000, // Color (5, 3, 2) (7, 1)
        8'b00001000, // Color (5, 3, 2) (8, 1)
        8'b00001000, // Color (5, 3, 2) (9, 1)
        8'b00000110, // Color (7, 5, 3) (10, 1)
        8'b00000110, // Color (7, 5, 3) (11, 1)
        8'b00001000, // Color (5, 3, 2) (12, 1)
        8'b00001000, // Color (5, 3, 2) (13, 1)
        8'b00001000, // Color (5, 3, 2) (14, 1)
        8'b01010110, // Color (2, 2, 2) (15, 1)
        8'b01010110, // Color (2, 2, 2) (0, 2)
        8'b00001000, // Color (5, 3, 2) (1, 2)
        8'b00000110, // Color (7, 5, 3) (2, 2)
        8'b01011000, // Color (9, 5, 4) (3, 2)
        8'b01011000, // Color (9, 5, 4) (4, 2)
        8'b01011000, // Color (9, 5, 4) (5, 2)
        8'b00000110, // Color (7, 5, 3) (6, 2)
        8'b00001000, // Color (5, 3, 2) (7, 2)
        8'b00001000, // Color (5, 3, 2) (8, 2)
        8'b00000110, // Color (7, 5, 3) (9, 2)
        8'b01011000, // Color (9, 5, 4) (10, 2)
        8'b01011000, // Color (9, 5, 4) (11, 2)
        8'b01011000, // Color (9, 5, 4) (12, 2)
        8'b00000110, // Color (7, 5, 3) (13, 2)
        8'b00001000, // Color (5, 3, 2) (14, 2)
        8'b01011110, // Color (3, 2, 2) (15, 2)
        8'b01011110, // Color (3, 2, 2) (0, 3)
        8'b00001000, // Color (5, 3, 2) (1, 3)
        8'b01011000, // Color (9, 5, 4) (2, 3)
        8'b00000110, // Color (7, 5, 3) (3, 3)
        8'b00000110, // Color (7, 5, 3) (4, 3)
        8'b00000110, // Color (7, 5, 3) (5, 3)
        8'b00001000, // Color (5, 3, 2) (6, 3)
        8'b01010110, // Color (2, 2, 2) (7, 3)
        8'b01010110, // Color (2, 2, 2) (8, 3)
        8'b00001000, // Color (5, 3, 2) (9, 3)
        8'b00000110, // Color (7, 5, 3) (10, 3)
        8'b00000110, // Color (7, 5, 3) (11, 3)
        8'b00000110, // Color (7, 5, 3) (12, 3)
        8'b01011000, // Color (9, 5, 4) (13, 3)
        8'b00001000, // Color (5, 3, 2) (14, 3)
        8'b01011110, // Color (3, 2, 2) (15, 3)
        8'b01011110, // Color (3, 2, 2) (0, 4)
        8'b00001000, // Color (5, 3, 2) (1, 4)
        8'b01011000, // Color (9, 5, 4) (2, 4)
        8'b00000110, // Color (7, 5, 3) (3, 4)
        8'b00000110, // Color (7, 5, 3) (4, 4)
        8'b00000110, // Color (7, 5, 3) (5, 4)
        8'b00001000, // Color (5, 3, 2) (6, 4)
        8'b01010110, // Color (2, 2, 2) (7, 4)
        8'b01100000, // Color (1, 1, 1) (8, 4)
        8'b00001000, // Color (5, 3, 2) (9, 4)
        8'b00000110, // Color (7, 5, 3) (10, 4)
        8'b00000110, // Color (7, 5, 3) (11, 4)
        8'b00000110, // Color (7, 5, 3) (12, 4)
        8'b01011000, // Color (9, 5, 4) (13, 4)
        8'b00000110, // Color (7, 5, 3) (14, 4)
        8'b01011110, // Color (3, 2, 2) (15, 4)
        8'b01010110, // Color (2, 2, 2) (0, 5)
        8'b00001000, // Color (5, 3, 2) (1, 5)
        8'b01011000, // Color (9, 5, 4) (2, 5)
        8'b00000110, // Color (7, 5, 3) (3, 5)
        8'b00000110, // Color (7, 5, 3) (4, 5)
        8'b00000110, // Color (7, 5, 3) (5, 5)
        8'b00001000, // Color (5, 3, 2) (6, 5)
        8'b01100000, // Color (1, 1, 1) (7, 5)
        8'b01100000, // Color (1, 1, 1) (8, 5)
        8'b00001000, // Color (5, 3, 2) (9, 5)
        8'b00000110, // Color (7, 5, 3) (10, 5)
        8'b00000110, // Color (7, 5, 3) (11, 5)
        8'b00000110, // Color (7, 5, 3) (12, 5)
        8'b01011000, // Color (9, 5, 4) (13, 5)
        8'b00000110, // Color (7, 5, 3) (14, 5)
        8'b01011110, // Color (3, 2, 2) (15, 5)
        8'b01010110, // Color (2, 2, 2) (0, 6)
        8'b00001000, // Color (5, 3, 2) (1, 6)
        8'b01011000, // Color (9, 5, 4) (2, 6)
        8'b00000110, // Color (7, 5, 3) (3, 6)
        8'b00000110, // Color (7, 5, 3) (4, 6)
        8'b00000110, // Color (7, 5, 3) (5, 6)
        8'b00001000, // Color (5, 3, 2) (6, 6)
        8'b01100000, // Color (1, 1, 1) (7, 6)
        8'b01100000, // Color (1, 1, 1) (8, 6)
        8'b00001000, // Color (5, 3, 2) (9, 6)
        8'b00000110, // Color (7, 5, 3) (10, 6)
        8'b00000110, // Color (7, 5, 3) (11, 6)
        8'b00000110, // Color (7, 5, 3) (12, 6)
        8'b01011000, // Color (9, 5, 4) (13, 6)
        8'b00000110, // Color (7, 5, 3) (14, 6)
        8'b01011110, // Color (3, 2, 2) (15, 6)
        8'b01011110, // Color (3, 2, 2) (0, 7)
        8'b00000110, // Color (7, 5, 3) (1, 7)
        8'b01011000, // Color (9, 5, 4) (2, 7)
        8'b00000110, // Color (7, 5, 3) (3, 7)
        8'b00000110, // Color (7, 5, 3) (4, 7)
        8'b00000110, // Color (7, 5, 3) (5, 7)
        8'b00001000, // Color (5, 3, 2) (6, 7)
        8'b01100000, // Color (1, 1, 1) (7, 7)
        8'b01100000, // Color (1, 1, 1) (8, 7)
        8'b00001000, // Color (5, 3, 2) (9, 7)
        8'b00000110, // Color (7, 5, 3) (10, 7)
        8'b00000110, // Color (7, 5, 3) (11, 7)
        8'b00000110, // Color (7, 5, 3) (12, 7)
        8'b01011000, // Color (9, 5, 4) (13, 7)
        8'b00001000, // Color (5, 3, 2) (14, 7)
        8'b01011110, // Color (3, 2, 2) (15, 7)
        8'b01011110, // Color (3, 2, 2) (0, 8)
        8'b00000110, // Color (7, 5, 3) (1, 8)
        8'b01011000, // Color (9, 5, 4) (2, 8)
        8'b00000110, // Color (7, 5, 3) (3, 8)
        8'b00000110, // Color (7, 5, 3) (4, 8)
        8'b00000110, // Color (7, 5, 3) (5, 8)
        8'b00001000, // Color (5, 3, 2) (6, 8)
        8'b01100000, // Color (1, 1, 1) (7, 8)
        8'b01100000, // Color (1, 1, 1) (8, 8)
        8'b00001000, // Color (5, 3, 2) (9, 8)
        8'b00000110, // Color (7, 5, 3) (10, 8)
        8'b00000110, // Color (7, 5, 3) (11, 8)
        8'b00000110, // Color (7, 5, 3) (12, 8)
        8'b01011000, // Color (9, 5, 4) (13, 8)
        8'b00001000, // Color (5, 3, 2) (14, 8)
        8'b01011110, // Color (3, 2, 2) (15, 8)
        8'b01011110, // Color (3, 2, 2) (0, 9)
        8'b00000110, // Color (7, 5, 3) (1, 9)
        8'b01011000, // Color (9, 5, 4) (2, 9)
        8'b00000110, // Color (7, 5, 3) (3, 9)
        8'b00000110, // Color (7, 5, 3) (4, 9)
        8'b00000110, // Color (7, 5, 3) (5, 9)
        8'b00001000, // Color (5, 3, 2) (6, 9)
        8'b01100000, // Color (1, 1, 1) (7, 9)
        8'b01100000, // Color (1, 1, 1) (8, 9)
        8'b00001000, // Color (5, 3, 2) (9, 9)
        8'b00000110, // Color (7, 5, 3) (10, 9)
        8'b00000110, // Color (7, 5, 3) (11, 9)
        8'b00000110, // Color (7, 5, 3) (12, 9)
        8'b01011000, // Color (9, 5, 4) (13, 9)
        8'b00001000, // Color (5, 3, 2) (14, 9)
        8'b01011110, // Color (3, 2, 2) (15, 9)
        8'b01011110, // Color (3, 2, 2) (0, 10)
        8'b00001000, // Color (5, 3, 2) (1, 10)
        8'b01011000, // Color (9, 5, 4) (2, 10)
        8'b00000110, // Color (7, 5, 3) (3, 10)
        8'b00000110, // Color (7, 5, 3) (4, 10)
        8'b00000110, // Color (7, 5, 3) (5, 10)
        8'b00001000, // Color (5, 3, 2) (6, 10)
        8'b01100000, // Color (1, 1, 1) (7, 10)
        8'b01100000, // Color (1, 1, 1) (8, 10)
        8'b00001000, // Color (5, 3, 2) (9, 10)
        8'b00000110, // Color (7, 5, 3) (10, 10)
        8'b00000110, // Color (7, 5, 3) (11, 10)
        8'b00000110, // Color (7, 5, 3) (12, 10)
        8'b01011000, // Color (9, 5, 4) (13, 10)
        8'b00000110, // Color (7, 5, 3) (14, 10)
        8'b01010110, // Color (2, 2, 2) (15, 10)
        8'b01011110, // Color (3, 2, 2) (0, 11)
        8'b00001000, // Color (5, 3, 2) (1, 11)
        8'b01011000, // Color (9, 5, 4) (2, 11)
        8'b00000110, // Color (7, 5, 3) (3, 11)
        8'b00000110, // Color (7, 5, 3) (4, 11)
        8'b00000110, // Color (7, 5, 3) (5, 11)
        8'b00001000, // Color (5, 3, 2) (6, 11)
        8'b01100000, // Color (1, 1, 1) (7, 11)
        8'b01010110, // Color (2, 2, 2) (8, 11)
        8'b00001000, // Color (5, 3, 2) (9, 11)
        8'b00000110, // Color (7, 5, 3) (10, 11)
        8'b00000110, // Color (7, 5, 3) (11, 11)
        8'b00000110, // Color (7, 5, 3) (12, 11)
        8'b01011000, // Color (9, 5, 4) (13, 11)
        8'b00000110, // Color (7, 5, 3) (14, 11)
        8'b01010110, // Color (2, 2, 2) (15, 11)
        8'b01011110, // Color (3, 2, 2) (0, 12)
        8'b00001000, // Color (5, 3, 2) (1, 12)
        8'b01011000, // Color (9, 5, 4) (2, 12)
        8'b00000110, // Color (7, 5, 3) (3, 12)
        8'b00000110, // Color (7, 5, 3) (4, 12)
        8'b00000110, // Color (7, 5, 3) (5, 12)
        8'b00001000, // Color (5, 3, 2) (6, 12)
        8'b01010110, // Color (2, 2, 2) (7, 12)
        8'b01010110, // Color (2, 2, 2) (8, 12)
        8'b00001000, // Color (5, 3, 2) (9, 12)
        8'b00000110, // Color (7, 5, 3) (10, 12)
        8'b00000110, // Color (7, 5, 3) (11, 12)
        8'b00000110, // Color (7, 5, 3) (12, 12)
        8'b01011000, // Color (9, 5, 4) (13, 12)
        8'b00000110, // Color (7, 5, 3) (14, 12)
        8'b01011110, // Color (3, 2, 2) (15, 12)
        8'b01011110, // Color (3, 2, 2) (0, 13)
        8'b00001000, // Color (5, 3, 2) (1, 13)
        8'b00000110, // Color (7, 5, 3) (2, 13)
        8'b01011000, // Color (9, 5, 4) (3, 13)
        8'b01011000, // Color (9, 5, 4) (4, 13)
        8'b01011000, // Color (9, 5, 4) (5, 13)
        8'b00000110, // Color (7, 5, 3) (6, 13)
        8'b00001000, // Color (5, 3, 2) (7, 13)
        8'b00001000, // Color (5, 3, 2) (8, 13)
        8'b00000110, // Color (7, 5, 3) (9, 13)
        8'b01011000, // Color (9, 5, 4) (10, 13)
        8'b01011000, // Color (9, 5, 4) (11, 13)
        8'b01011000, // Color (9, 5, 4) (12, 13)
        8'b00000110, // Color (7, 5, 3) (13, 13)
        8'b00001000, // Color (5, 3, 2) (14, 13)
        8'b01011110, // Color (3, 2, 2) (15, 13)
        8'b01010110, // Color (2, 2, 2) (0, 14)
        8'b00001000, // Color (5, 3, 2) (1, 14)
        8'b00001000, // Color (5, 3, 2) (2, 14)
        8'b00000110, // Color (7, 5, 3) (3, 14)
        8'b00000110, // Color (7, 5, 3) (4, 14)
        8'b00001000, // Color (5, 3, 2) (5, 14)
        8'b00001000, // Color (5, 3, 2) (6, 14)
        8'b00001000, // Color (5, 3, 2) (7, 14)
        8'b00000110, // Color (7, 5, 3) (8, 14)
        8'b00000110, // Color (7, 5, 3) (9, 14)
        8'b00000110, // Color (7, 5, 3) (10, 14)
        8'b00001000, // Color (5, 3, 2) (11, 14)
        8'b00001000, // Color (5, 3, 2) (12, 14)
        8'b00001000, // Color (5, 3, 2) (13, 14)
        8'b00001000, // Color (5, 3, 2) (14, 14)
        8'b01010110, // Color (2, 2, 2) (15, 14)
        8'b01010110, // Color (2, 2, 2) (0, 15)
        8'b01010110, // Color (2, 2, 2) (1, 15)
        8'b01010110, // Color (2, 2, 2) (2, 15)
        8'b01011110, // Color (3, 2, 2) (3, 15)
        8'b01011110, // Color (3, 2, 2) (4, 15)
        8'b01011110, // Color (3, 2, 2) (5, 15)
        8'b01011110, // Color (3, 2, 2) (6, 15)
        8'b01011110, // Color (3, 2, 2) (7, 15)
        8'b01011110, // Color (3, 2, 2) (8, 15)
        8'b01011110, // Color (3, 2, 2) (9, 15)
        8'b01011110, // Color (3, 2, 2) (10, 15)
        8'b01010110, // Color (2, 2, 2) (11, 15)
        8'b01011110, // Color (3, 2, 2) (12, 15)
        8'b01010110, // Color (2, 2, 2) (13, 15)
        8'b01010110, // Color (2, 2, 2) (14, 15)
        8'b01010110, // Color (2, 2, 2) (15, 15)
        // 10_cobblestone
        8'b00001100, // Color (6, 6, 6) (0, 0)
        8'b00001100, // Color (6, 6, 6) (1, 0)
        8'b01100010, // Color (10, 10, 10) (2, 0)
        8'b01100010, // Color (10, 10, 10) (3, 0)
        8'b01100100, // Color (5, 5, 5) (4, 0)
        8'b00001100, // Color (6, 6, 6) (5, 0)
        8'b00001100, // Color (6, 6, 6) (6, 0)
        8'b01100010, // Color (10, 10, 10) (7, 0)
        8'b01100110, // Color (11, 11, 11) (8, 0)
        8'b01100010, // Color (10, 10, 10) (9, 0)
        8'b00001010, // Color (8, 8, 8) (10, 0)
        8'b00001100, // Color (6, 6, 6) (11, 0)
        8'b00001010, // Color (8, 8, 8) (12, 0)
        8'b01100110, // Color (11, 11, 11) (13, 0)
        8'b01100010, // Color (10, 10, 10) (14, 0)
        8'b00001010, // Color (8, 8, 8) (15, 0)
        8'b00001100, // Color (6, 6, 6) (0, 1)
        8'b01100010, // Color (10, 10, 10) (1, 1)
        8'b01100110, // Color (11, 11, 11) (2, 1)
        8'b00001010, // Color (8, 8, 8) (3, 1)
        8'b00001010, // Color (8, 8, 8) (4, 1)
        8'b01100100, // Color (5, 5, 5) (5, 1)
        8'b01100110, // Color (11, 11, 11) (6, 1)
        8'b01100110, // Color (11, 11, 11) (7, 1)
        8'b01100010, // Color (10, 10, 10) (8, 1)
        8'b00001010, // Color (8, 8, 8) (9, 1)
        8'b00001010, // Color (8, 8, 8) (10, 1)
        8'b01100100, // Color (5, 5, 5) (11, 1)
        8'b00001100, // Color (6, 6, 6) (12, 1)
        8'b00001010, // Color (8, 8, 8) (13, 1)
        8'b00001100, // Color (6, 6, 6) (14, 1)
        8'b00001010, // Color (8, 8, 8) (15, 1)
        8'b00001100, // Color (6, 6, 6) (0, 2)
        8'b01100010, // Color (10, 10, 10) (1, 2)
        8'b00001010, // Color (8, 8, 8) (2, 2)
        8'b01100010, // Color (10, 10, 10) (3, 2)
        8'b00001100, // Color (6, 6, 6) (4, 2)
        8'b00001100, // Color (6, 6, 6) (5, 2)
        8'b01100010, // Color (10, 10, 10) (6, 2)
        8'b00001010, // Color (8, 8, 8) (7, 2)
        8'b00001010, // Color (8, 8, 8) (8, 2)
        8'b01100010, // Color (10, 10, 10) (9, 2)
        8'b00001100, // Color (6, 6, 6) (10, 2)
        8'b00001100, // Color (6, 6, 6) (11, 2)
        8'b01100100, // Color (5, 5, 5) (12, 2)
        8'b00001100, // Color (6, 6, 6) (13, 2)
        8'b00001010, // Color (8, 8, 8) (14, 2)
        8'b00001100, // Color (6, 6, 6) (15, 2)
        8'b00001100, // Color (6, 6, 6) (0, 3)
        8'b00001100, // Color (6, 6, 6) (1, 3)
        8'b00001010, // Color (8, 8, 8) (2, 3)
        8'b00001100, // Color (6, 6, 6) (3, 3)
        8'b00001100, // Color (6, 6, 6) (4, 3)
        8'b00001100, // Color (6, 6, 6) (5, 3)
        8'b00001010, // Color (8, 8, 8) (6, 3)
        8'b00001100, // Color (6, 6, 6) (7, 3)
        8'b00001010, // Color (8, 8, 8) (8, 3)
        8'b00001100, // Color (6, 6, 6) (9, 3)
        8'b00001100, // Color (6, 6, 6) (10, 3)
        8'b00001010, // Color (8, 8, 8) (11, 3)
        8'b01100010, // Color (10, 10, 10) (12, 3)
        8'b00001010, // Color (8, 8, 8) (13, 3)
        8'b00001100, // Color (6, 6, 6) (14, 3)
        8'b01100100, // Color (5, 5, 5) (15, 3)
        8'b01100100, // Color (5, 5, 5) (0, 4)
        8'b00001100, // Color (6, 6, 6) (1, 4)
        8'b00001100, // Color (6, 6, 6) (2, 4)
        8'b00001010, // Color (8, 8, 8) (3, 4)
        8'b01100110, // Color (11, 11, 11) (4, 4)
        8'b01100010, // Color (10, 10, 10) (5, 4)
        8'b00001100, // Color (6, 6, 6) (6, 4)
        8'b00001010, // Color (8, 8, 8) (7, 4)
        8'b00001100, // Color (6, 6, 6) (8, 4)
        8'b00001100, // Color (6, 6, 6) (9, 4)
        8'b01100110, // Color (11, 11, 11) (10, 4)
        8'b01100010, // Color (10, 10, 10) (11, 4)
        8'b01100010, // Color (10, 10, 10) (12, 4)
        8'b01100010, // Color (10, 10, 10) (13, 4)
        8'b00001010, // Color (8, 8, 8) (14, 4)
        8'b00001100, // Color (6, 6, 6) (15, 4)
        8'b01100110, // Color (11, 11, 11) (0, 5)
        8'b00001100, // Color (6, 6, 6) (1, 5)
        8'b01100010, // Color (10, 10, 10) (2, 5)
        8'b01100110, // Color (11, 11, 11) (3, 5)
        8'b00001010, // Color (8, 8, 8) (4, 5)
        8'b00001010, // Color (8, 8, 8) (5, 5)
        8'b00001100, // Color (6, 6, 6) (6, 5)
        8'b00001100, // Color (6, 6, 6) (7, 5)
        8'b01100100, // Color (5, 5, 5) (8, 5)
        8'b00001010, // Color (8, 8, 8) (9, 5)
        8'b00001010, // Color (8, 8, 8) (10, 5)
        8'b01100110, // Color (11, 11, 11) (11, 5)
        8'b01100010, // Color (10, 10, 10) (12, 5)
        8'b00001010, // Color (8, 8, 8) (13, 5)
        8'b00001100, // Color (6, 6, 6) (14, 5)
        8'b00001010, // Color (8, 8, 8) (15, 5)
        8'b01100010, // Color (10, 10, 10) (0, 6)
        8'b00001010, // Color (8, 8, 8) (1, 6)
        8'b00001100, // Color (6, 6, 6) (2, 6)
        8'b00001010, // Color (8, 8, 8) (3, 6)
        8'b01100010, // Color (10, 10, 10) (4, 6)
        8'b00001010, // Color (8, 8, 8) (5, 6)
        8'b00001010, // Color (8, 8, 8) (6, 6)
        8'b00001100, // Color (6, 6, 6) (7, 6)
        8'b00001100, // Color (6, 6, 6) (8, 6)
        8'b00001100, // Color (6, 6, 6) (9, 6)
        8'b00001100, // Color (6, 6, 6) (10, 6)
        8'b01100010, // Color (10, 10, 10) (11, 6)
        8'b00001010, // Color (8, 8, 8) (12, 6)
        8'b00001100, // Color (6, 6, 6) (13, 6)
        8'b00001100, // Color (6, 6, 6) (14, 6)
        8'b01100110, // Color (11, 11, 11) (15, 6)
        8'b00001010, // Color (8, 8, 8) (0, 7)
        8'b00001010, // Color (8, 8, 8) (1, 7)
        8'b00001100, // Color (6, 6, 6) (2, 7)
        8'b00001100, // Color (6, 6, 6) (3, 7)
        8'b00001010, // Color (8, 8, 8) (4, 7)
        8'b00001010, // Color (8, 8, 8) (5, 7)
        8'b00001100, // Color (6, 6, 6) (6, 7)
        8'b00001100, // Color (6, 6, 6) (7, 7)
        8'b00001010, // Color (8, 8, 8) (8, 7)
        8'b01100110, // Color (11, 11, 11) (9, 7)
        8'b01100010, // Color (10, 10, 10) (10, 7)
        8'b00001100, // Color (6, 6, 6) (11, 7)
        8'b00001100, // Color (6, 6, 6) (12, 7)
        8'b00001010, // Color (8, 8, 8) (13, 7)
        8'b00001100, // Color (6, 6, 6) (14, 7)
        8'b00001010, // Color (8, 8, 8) (15, 7)
        8'b00001100, // Color (6, 6, 6) (0, 8)
        8'b00001100, // Color (6, 6, 6) (1, 8)
        8'b01100110, // Color (11, 11, 11) (2, 8)
        8'b01100010, // Color (10, 10, 10) (3, 8)
        8'b00001100, // Color (6, 6, 6) (4, 8)
        8'b00001100, // Color (6, 6, 6) (5, 8)
        8'b00001100, // Color (6, 6, 6) (6, 8)
        8'b00001010, // Color (8, 8, 8) (7, 8)
        8'b01100110, // Color (11, 11, 11) (8, 8)
        8'b00001010, // Color (8, 8, 8) (9, 8)
        8'b00001010, // Color (8, 8, 8) (10, 8)
        8'b00001010, // Color (8, 8, 8) (11, 8)
        8'b00001100, // Color (6, 6, 6) (12, 8)
        8'b00001100, // Color (6, 6, 6) (13, 8)
        8'b01100100, // Color (5, 5, 5) (14, 8)
        8'b00001100, // Color (6, 6, 6) (15, 8)
        8'b00001100, // Color (6, 6, 6) (0, 9)
        8'b01100110, // Color (11, 11, 11) (1, 9)
        8'b01100010, // Color (10, 10, 10) (2, 9)
        8'b00001010, // Color (8, 8, 8) (3, 9)
        8'b00001100, // Color (6, 6, 6) (4, 9)
        8'b00001010, // Color (8, 8, 8) (5, 9)
        8'b00001100, // Color (6, 6, 6) (6, 9)
        8'b00001100, // Color (6, 6, 6) (7, 9)
        8'b00001010, // Color (8, 8, 8) (8, 9)
        8'b00001010, // Color (8, 8, 8) (9, 9)
        8'b00001100, // Color (6, 6, 6) (10, 9)
        8'b00001100, // Color (6, 6, 6) (11, 9)
        8'b00001100, // Color (6, 6, 6) (12, 9)
        8'b00001010, // Color (8, 8, 8) (13, 9)
        8'b01100010, // Color (10, 10, 10) (14, 9)
        8'b00001100, // Color (6, 6, 6) (15, 9)
        8'b00001010, // Color (8, 8, 8) (0, 10)
        8'b00001100, // Color (6, 6, 6) (1, 10)
        8'b00001010, // Color (8, 8, 8) (2, 10)
        8'b00001100, // Color (6, 6, 6) (3, 10)
        8'b00001010, // Color (8, 8, 8) (4, 10)
        8'b00001100, // Color (6, 6, 6) (5, 10)
        8'b00001100, // Color (6, 6, 6) (6, 10)
        8'b01100100, // Color (5, 5, 5) (7, 10)
        8'b00001100, // Color (6, 6, 6) (8, 10)
        8'b00001100, // Color (6, 6, 6) (9, 10)
        8'b00001100, // Color (6, 6, 6) (10, 10)
        8'b00001100, // Color (6, 6, 6) (11, 10)
        8'b01100100, // Color (5, 5, 5) (12, 10)
        8'b01100010, // Color (10, 10, 10) (13, 10)
        8'b01100010, // Color (10, 10, 10) (14, 10)
        8'b01100110, // Color (11, 11, 11) (15, 10)
        8'b00001010, // Color (8, 8, 8) (0, 11)
        8'b00001100, // Color (6, 6, 6) (1, 11)
        8'b00001100, // Color (6, 6, 6) (2, 11)
        8'b00001100, // Color (6, 6, 6) (3, 11)
        8'b00001100, // Color (6, 6, 6) (4, 11)
        8'b00001100, // Color (6, 6, 6) (5, 11)
        8'b00001010, // Color (8, 8, 8) (6, 11)
        8'b01100110, // Color (11, 11, 11) (7, 11)
        8'b01100010, // Color (10, 10, 10) (8, 11)
        8'b00001100, // Color (6, 6, 6) (9, 11)
        8'b00001100, // Color (6, 6, 6) (10, 11)
        8'b01100100, // Color (5, 5, 5) (11, 11)
        8'b00001010, // Color (8, 8, 8) (12, 11)
        8'b01100110, // Color (11, 11, 11) (13, 11)
        8'b01100110, // Color (11, 11, 11) (14, 11)
        8'b00001010, // Color (8, 8, 8) (15, 11)
        8'b00001100, // Color (6, 6, 6) (0, 12)
        8'b00001010, // Color (8, 8, 8) (1, 12)
        8'b01100110, // Color (11, 11, 11) (2, 12)
        8'b01100010, // Color (10, 10, 10) (3, 12)
        8'b00001100, // Color (6, 6, 6) (4, 12)
        8'b00001100, // Color (6, 6, 6) (5, 12)
        8'b01100110, // Color (11, 11, 11) (6, 12)
        8'b01100010, // Color (10, 10, 10) (7, 12)
        8'b00001010, // Color (8, 8, 8) (8, 12)
        8'b01100010, // Color (10, 10, 10) (9, 12)
        8'b00001100, // Color (6, 6, 6) (10, 12)
        8'b00001100, // Color (6, 6, 6) (11, 12)
        8'b00001010, // Color (8, 8, 8) (12, 12)
        8'b00001010, // Color (8, 8, 8) (13, 12)
        8'b00001100, // Color (6, 6, 6) (14, 12)
        8'b00001010, // Color (8, 8, 8) (15, 12)
        8'b00001100, // Color (6, 6, 6) (0, 13)
        8'b01100110, // Color (11, 11, 11) (1, 13)
        8'b01100010, // Color (10, 10, 10) (2, 13)
        8'b00001010, // Color (8, 8, 8) (3, 13)
        8'b00001010, // Color (8, 8, 8) (4, 13)
        8'b00001100, // Color (6, 6, 6) (5, 13)
        8'b01100010, // Color (10, 10, 10) (6, 13)
        8'b00001010, // Color (8, 8, 8) (7, 13)
        8'b00001100, // Color (6, 6, 6) (8, 13)
        8'b00001010, // Color (8, 8, 8) (9, 13)
        8'b00001010, // Color (8, 8, 8) (10, 13)
        8'b00001100, // Color (6, 6, 6) (11, 13)
        8'b00001100, // Color (6, 6, 6) (12, 13)
        8'b00001100, // Color (6, 6, 6) (13, 13)
        8'b00001010, // Color (8, 8, 8) (14, 13)
        8'b00001100, // Color (6, 6, 6) (15, 13)
        8'b01100010, // Color (10, 10, 10) (0, 14)
        8'b01100010, // Color (10, 10, 10) (1, 14)
        8'b00001010, // Color (8, 8, 8) (2, 14)
        8'b00001100, // Color (6, 6, 6) (3, 14)
        8'b00001010, // Color (8, 8, 8) (4, 14)
        8'b00001100, // Color (6, 6, 6) (5, 14)
        8'b00001100, // Color (6, 6, 6) (6, 14)
        8'b00001100, // Color (6, 6, 6) (7, 14)
        8'b00001010, // Color (8, 8, 8) (8, 14)
        8'b00001010, // Color (8, 8, 8) (9, 14)
        8'b00001100, // Color (6, 6, 6) (10, 14)
        8'b00001100, // Color (6, 6, 6) (11, 14)
        8'b01100010, // Color (10, 10, 10) (12, 14)
        8'b00001010, // Color (8, 8, 8) (13, 14)
        8'b00001100, // Color (6, 6, 6) (14, 14)
        8'b00001100, // Color (6, 6, 6) (15, 14)
        8'b00001100, // Color (6, 6, 6) (0, 15)
        8'b00001010, // Color (8, 8, 8) (1, 15)
        8'b00001100, // Color (6, 6, 6) (2, 15)
        8'b00001100, // Color (6, 6, 6) (3, 15)
        8'b00001100, // Color (6, 6, 6) (4, 15)
        8'b00001010, // Color (8, 8, 8) (5, 15)
        8'b00001100, // Color (6, 6, 6) (6, 15)
        8'b00001100, // Color (6, 6, 6) (7, 15)
        8'b00001100, // Color (6, 6, 6) (8, 15)
        8'b00001100, // Color (6, 6, 6) (9, 15)
        8'b00001100, // Color (6, 6, 6) (10, 15)
        8'b00001010, // Color (8, 8, 8) (11, 15)
        8'b01100110, // Color (11, 11, 11) (12, 15)
        8'b01100010, // Color (10, 10, 10) (13, 15)
        8'b00001010, // Color (8, 8, 8) (14, 15)
        8'b00001100, // Color (6, 6, 6) (15, 15)
        // 11_crafting_table_front
        8'b01101000, // Color (1, 1, 0) (0, 0)
        8'b00111100, // Color (10, 8, 5) (1, 0)
        8'b00111010, // Color (11, 9, 5) (2, 0)
        8'b00111110, // Color (12, 9, 6) (3, 0)
        8'b00111110, // Color (12, 9, 6) (4, 0)
        8'b00110110, // Color (3, 2, 1) (5, 0)
        8'b01101010, // Color (7, 3, 2) (6, 0)
        8'b01011010, // Color (4, 2, 1) (7, 0)
        8'b01011010, // Color (4, 2, 1) (8, 0)
        8'b01101010, // Color (7, 3, 2) (9, 0)
        8'b00110110, // Color (3, 2, 1) (10, 0)
        8'b00111110, // Color (12, 9, 6) (11, 0)
        8'b00111110, // Color (12, 9, 6) (12, 0)
        8'b00111110, // Color (12, 9, 6) (13, 0)
        8'b00111010, // Color (11, 9, 5) (14, 0)
        8'b01101000, // Color (1, 1, 0) (15, 0)
        8'b01101000, // Color (1, 1, 0) (0, 1)
        8'b00111010, // Color (11, 9, 5) (1, 1)
        8'b00111100, // Color (10, 8, 5) (2, 1)
        8'b00111100, // Color (10, 8, 5) (3, 1)
        8'b00110100, // Color (9, 7, 4) (4, 1)
        8'b01000010, // Color (9, 8, 4) (5, 1)
        8'b00110110, // Color (3, 2, 1) (6, 1)
        8'b01011010, // Color (4, 2, 1) (7, 1)
        8'b01011010, // Color (4, 2, 1) (8, 1)
        8'b00110110, // Color (3, 2, 1) (9, 1)
        8'b00111100, // Color (10, 8, 5) (10, 1)
        8'b00111100, // Color (10, 8, 5) (11, 1)
        8'b00111010, // Color (11, 9, 5) (12, 1)
        8'b00111010, // Color (11, 9, 5) (13, 1)
        8'b01000010, // Color (9, 8, 4) (14, 1)
        8'b01101000, // Color (1, 1, 0) (15, 1)
        8'b01101000, // Color (1, 1, 0) (0, 2)
        8'b00111010, // Color (11, 9, 5) (1, 2)
        8'b00111010, // Color (11, 9, 5) (2, 2)
        8'b00111010, // Color (11, 9, 5) (3, 2)
        8'b00111100, // Color (10, 8, 5) (4, 2)
        8'b00111010, // Color (11, 9, 5) (5, 2)
        8'b00111100, // Color (10, 8, 5) (6, 2)
        8'b00110110, // Color (3, 2, 1) (7, 2)
        8'b00110110, // Color (3, 2, 1) (8, 2)
        8'b01000010, // Color (9, 8, 4) (9, 2)
        8'b01000010, // Color (9, 8, 4) (10, 2)
        8'b00111100, // Color (10, 8, 5) (11, 2)
        8'b00111100, // Color (10, 8, 5) (12, 2)
        8'b00111010, // Color (11, 9, 5) (13, 2)
        8'b00111010, // Color (11, 9, 5) (14, 2)
        8'b01101000, // Color (1, 1, 0) (15, 2)
        8'b01101000, // Color (1, 1, 0) (0, 3)
        8'b01000000, // Color (7, 6, 3) (1, 3)
        8'b01000000, // Color (7, 6, 3) (2, 3)
        8'b00110100, // Color (9, 7, 4) (3, 3)
        8'b00110100, // Color (9, 7, 4) (4, 3)
        8'b01000000, // Color (7, 6, 3) (5, 3)
        8'b01000100, // Color (6, 5, 2) (6, 3)
        8'b01101000, // Color (1, 1, 0) (7, 3)
        8'b01101000, // Color (1, 1, 0) (8, 3)
        8'b01000000, // Color (7, 6, 3) (9, 3)
        8'b01000100, // Color (6, 5, 2) (10, 3)
        8'b01101100, // Color (4, 2, 0) (11, 3)
        8'b01101100, // Color (4, 2, 0) (12, 3)
        8'b01101100, // Color (4, 2, 0) (13, 3)
        8'b01000000, // Color (7, 6, 3) (14, 3)
        8'b01101000, // Color (1, 1, 0) (15, 3)
        8'b01101000, // Color (1, 1, 0) (0, 4)
        8'b00111110, // Color (12, 9, 6) (1, 4)
        8'b01000010, // Color (9, 8, 4) (2, 4)
        8'b00111110, // Color (12, 9, 6) (3, 4)
        8'b00111110, // Color (12, 9, 6) (4, 4)
        8'b00111110, // Color (12, 9, 6) (5, 4)
        8'b00111110, // Color (12, 9, 6) (6, 4)
        8'b01011010, // Color (4, 2, 1) (7, 4)
        8'b01011010, // Color (4, 2, 1) (8, 4)
        8'b00111110, // Color (12, 9, 6) (9, 4)
        8'b00111110, // Color (12, 9, 6) (10, 4)
        8'b01101110, // Color (2, 1, 0) (11, 4)
        8'b00111100, // Color (10, 8, 5) (12, 4)
        8'b01101110, // Color (2, 1, 0) (13, 4)
        8'b01000010, // Color (9, 8, 4) (14, 4)
        8'b01101000, // Color (1, 1, 0) (15, 4)
        8'b01101000, // Color (1, 1, 0) (0, 5)
        8'b00111010, // Color (11, 9, 5) (1, 5)
        8'b00111010, // Color (11, 9, 5) (2, 5)
        8'b01101100, // Color (4, 2, 0) (3, 5)
        8'b01000010, // Color (9, 8, 4) (4, 5)
        8'b00111100, // Color (10, 8, 5) (5, 5)
        8'b01000010, // Color (9, 8, 4) (6, 5)
        8'b00110110, // Color (3, 2, 1) (7, 5)
        8'b00110110, // Color (3, 2, 1) (8, 5)
        8'b00111100, // Color (10, 8, 5) (9, 5)
        8'b00111100, // Color (10, 8, 5) (10, 5)
        8'b01101110, // Color (2, 1, 0) (11, 5)
        8'b01101110, // Color (2, 1, 0) (12, 5)
        8'b01101110, // Color (2, 1, 0) (13, 5)
        8'b00111010, // Color (11, 9, 5) (14, 5)
        8'b01101000, // Color (1, 1, 0) (15, 5)
        8'b01101000, // Color (1, 1, 0) (0, 6)
        8'b01000010, // Color (9, 8, 4) (1, 6)
        8'b00111100, // Color (10, 8, 5) (2, 6)
        8'b01101110, // Color (2, 1, 0) (3, 6)
        8'b00111100, // Color (10, 8, 5) (4, 6)
        8'b00111100, // Color (10, 8, 5) (5, 6)
        8'b00111100, // Color (10, 8, 5) (6, 6)
        8'b00110110, // Color (3, 2, 1) (7, 6)
        8'b00110110, // Color (3, 2, 1) (8, 6)
        8'b00111010, // Color (11, 9, 5) (9, 6)
        8'b00111010, // Color (11, 9, 5) (10, 6)
        8'b01100110, // Color (11, 11, 11) (11, 6)
        8'b01100110, // Color (11, 11, 11) (12, 6)
        8'b01100110, // Color (11, 11, 11) (13, 6)
        8'b01000010, // Color (9, 8, 4) (14, 6)
        8'b01101000, // Color (1, 1, 0) (15, 6)
        8'b01101000, // Color (1, 1, 0) (0, 7)
        8'b01000100, // Color (6, 5, 2) (1, 7)
        8'b01000000, // Color (7, 6, 3) (2, 7)
        8'b01101110, // Color (2, 1, 0) (3, 7)
        8'b00110100, // Color (9, 7, 4) (4, 7)
        8'b01000000, // Color (7, 6, 3) (5, 7)
        8'b01000100, // Color (6, 5, 2) (6, 7)
        8'b01101000, // Color (1, 1, 0) (7, 7)
        8'b01101000, // Color (1, 1, 0) (8, 7)
        8'b01000100, // Color (6, 5, 2) (9, 7)
        8'b01000000, // Color (7, 6, 3) (10, 7)
        8'b01110000, // Color (15, 15, 15) (11, 7)
        8'b01110010, // Color (13, 13, 13) (12, 7)
        8'b01110010, // Color (13, 13, 13) (13, 7)
        8'b01000000, // Color (7, 6, 3) (14, 7)
        8'b01101000, // Color (1, 1, 0) (15, 7)
        8'b01101000, // Color (1, 1, 0) (0, 8)
        8'b00111110, // Color (12, 9, 6) (1, 8)
        8'b00111110, // Color (12, 9, 6) (2, 8)
        8'b01101110, // Color (2, 1, 0) (3, 8)
        8'b00111100, // Color (10, 8, 5) (4, 8)
        8'b00111100, // Color (10, 8, 5) (5, 8)
        8'b00111110, // Color (12, 9, 6) (6, 8)
        8'b01011010, // Color (4, 2, 1) (7, 8)
        8'b01011010, // Color (4, 2, 1) (8, 8)
        8'b00111110, // Color (12, 9, 6) (9, 8)
        8'b00111110, // Color (12, 9, 6) (10, 8)
        8'b01110000, // Color (15, 15, 15) (11, 8)
        8'b01110010, // Color (13, 13, 13) (12, 8)
        8'b01110010, // Color (13, 13, 13) (13, 8)
        8'b00111010, // Color (11, 9, 5) (14, 8)
        8'b01101000, // Color (1, 1, 0) (15, 8)
        8'b01101000, // Color (1, 1, 0) (0, 9)
        8'b00111100, // Color (10, 8, 5) (1, 9)
        8'b01110010, // Color (13, 13, 13) (2, 9)
        8'b01110010, // Color (13, 13, 13) (3, 9)
        8'b01110010, // Color (13, 13, 13) (4, 9)
        8'b00111010, // Color (11, 9, 5) (5, 9)
        8'b00111100, // Color (10, 8, 5) (6, 9)
        8'b00110110, // Color (3, 2, 1) (7, 9)
        8'b00110110, // Color (3, 2, 1) (8, 9)
        8'b01000010, // Color (9, 8, 4) (9, 9)
        8'b00111100, // Color (10, 8, 5) (10, 9)
        8'b01000010, // Color (9, 8, 4) (11, 9)
        8'b01110010, // Color (13, 13, 13) (12, 9)
        8'b01110010, // Color (13, 13, 13) (13, 9)
        8'b01000010, // Color (9, 8, 4) (14, 9)
        8'b01101000, // Color (1, 1, 0) (15, 9)
        8'b01101000, // Color (1, 1, 0) (0, 10)
        8'b00111010, // Color (11, 9, 5) (1, 10)
        8'b01100110, // Color (11, 11, 11) (2, 10)
        8'b01110010, // Color (13, 13, 13) (3, 10)
        8'b01110000, // Color (15, 15, 15) (4, 10)
        8'b01000010, // Color (9, 8, 4) (5, 10)
        8'b01000010, // Color (9, 8, 4) (6, 10)
        8'b00110110, // Color (3, 2, 1) (7, 10)
        8'b00110110, // Color (3, 2, 1) (8, 10)
        8'b00111100, // Color (10, 8, 5) (9, 10)
        8'b00111100, // Color (10, 8, 5) (10, 10)
        8'b00111100, // Color (10, 8, 5) (11, 10)
        8'b01110000, // Color (15, 15, 15) (12, 10)
        8'b01110010, // Color (13, 13, 13) (13, 10)
        8'b00111010, // Color (11, 9, 5) (14, 10)
        8'b01101000, // Color (1, 1, 0) (15, 10)
        8'b01101000, // Color (1, 1, 0) (0, 11)
        8'b01000100, // Color (6, 5, 2) (1, 11)
        8'b01000000, // Color (7, 6, 3) (2, 11)
        8'b00110100, // Color (9, 7, 4) (3, 11)
        8'b00110100, // Color (9, 7, 4) (4, 11)
        8'b01000000, // Color (7, 6, 3) (5, 11)
        8'b01000100, // Color (6, 5, 2) (6, 11)
        8'b01110100, // Color (1, 0, 0) (7, 11)
        8'b01110100, // Color (1, 0, 0) (8, 11)
        8'b01000000, // Color (7, 6, 3) (9, 11)
        8'b00110100, // Color (9, 7, 4) (10, 11)
        8'b01000000, // Color (7, 6, 3) (11, 11)
        8'b01000000, // Color (7, 6, 3) (12, 11)
        8'b01110010, // Color (13, 13, 13) (13, 11)
        8'b01000100, // Color (6, 5, 2) (14, 11)
        8'b01101000, // Color (1, 1, 0) (15, 11)
        8'b01101000, // Color (1, 1, 0) (0, 12)
        8'b01000010, // Color (9, 8, 4) (1, 12)
        8'b00111010, // Color (11, 9, 5) (2, 12)
        8'b00111110, // Color (12, 9, 6) (3, 12)
        8'b00111110, // Color (12, 9, 6) (4, 12)
        8'b00111010, // Color (11, 9, 5) (5, 12)
        8'b00111010, // Color (11, 9, 5) (6, 12)
        8'b01011010, // Color (4, 2, 1) (7, 12)
        8'b01011010, // Color (4, 2, 1) (8, 12)
        8'b00111110, // Color (12, 9, 6) (9, 12)
        8'b00111110, // Color (12, 9, 6) (10, 12)
        8'b01000010, // Color (9, 8, 4) (11, 12)
        8'b00111110, // Color (12, 9, 6) (12, 12)
        8'b01110000, // Color (15, 15, 15) (13, 12)
        8'b00111110, // Color (12, 9, 6) (14, 12)
        8'b01101000, // Color (1, 1, 0) (15, 12)
        8'b01101000, // Color (1, 1, 0) (0, 13)
        8'b00111100, // Color (10, 8, 5) (1, 13)
        8'b00111010, // Color (11, 9, 5) (2, 13)
        8'b00111010, // Color (11, 9, 5) (3, 13)
        8'b01000010, // Color (9, 8, 4) (4, 13)
        8'b01000010, // Color (9, 8, 4) (5, 13)
        8'b00111100, // Color (10, 8, 5) (6, 13)
        8'b00110110, // Color (3, 2, 1) (7, 13)
        8'b00110110, // Color (3, 2, 1) (8, 13)
        8'b00111010, // Color (11, 9, 5) (9, 13)
        8'b00111010, // Color (11, 9, 5) (10, 13)
        8'b00111100, // Color (10, 8, 5) (11, 13)
        8'b00111010, // Color (11, 9, 5) (12, 13)
        8'b00111100, // Color (10, 8, 5) (13, 13)
        8'b00111100, // Color (10, 8, 5) (14, 13)
        8'b01101000, // Color (1, 1, 0) (15, 13)
        8'b01101000, // Color (1, 1, 0) (0, 14)
        8'b01000010, // Color (9, 8, 4) (1, 14)
        8'b01000010, // Color (9, 8, 4) (2, 14)
        8'b00111100, // Color (10, 8, 5) (3, 14)
        8'b00111010, // Color (11, 9, 5) (4, 14)
        8'b00111100, // Color (10, 8, 5) (5, 14)
        8'b01000010, // Color (9, 8, 4) (6, 14)
        8'b00110110, // Color (3, 2, 1) (7, 14)
        8'b00110110, // Color (3, 2, 1) (8, 14)
        8'b00111010, // Color (11, 9, 5) (9, 14)
        8'b00111100, // Color (10, 8, 5) (10, 14)
        8'b01000010, // Color (9, 8, 4) (11, 14)
        8'b01000010, // Color (9, 8, 4) (12, 14)
        8'b01000010, // Color (9, 8, 4) (13, 14)
        8'b01000010, // Color (9, 8, 4) (14, 14)
        8'b01101000, // Color (1, 1, 0) (15, 14)
        8'b01101000, // Color (1, 1, 0) (0, 15)
        8'b01000000, // Color (7, 6, 3) (1, 15)
        8'b01000000, // Color (7, 6, 3) (2, 15)
        8'b01000100, // Color (6, 5, 2) (3, 15)
        8'b01000100, // Color (6, 5, 2) (4, 15)
        8'b01000000, // Color (7, 6, 3) (5, 15)
        8'b00110100, // Color (9, 7, 4) (6, 15)
        8'b01101000, // Color (1, 1, 0) (7, 15)
        8'b01101000, // Color (1, 1, 0) (8, 15)
        8'b01000000, // Color (7, 6, 3) (9, 15)
        8'b01000100, // Color (6, 5, 2) (10, 15)
        8'b01000000, // Color (7, 6, 3) (11, 15)
        8'b01000100, // Color (6, 5, 2) (12, 15)
        8'b01000100, // Color (6, 5, 2) (13, 15)
        8'b01000100, // Color (6, 5, 2) (14, 15)
        8'b01101000, // Color (1, 1, 0) (15, 15)
        // 12_crafting_table_side
        8'b01101000, // Color (1, 1, 0) (0, 0)
        8'b00111100, // Color (10, 8, 5) (1, 0)
        8'b00111010, // Color (11, 9, 5) (2, 0)
        8'b00111110, // Color (12, 9, 6) (3, 0)
        8'b00111110, // Color (12, 9, 6) (4, 0)
        8'b00110110, // Color (3, 2, 1) (5, 0)
        8'b01101010, // Color (7, 3, 2) (6, 0)
        8'b01011010, // Color (4, 2, 1) (7, 0)
        8'b01011010, // Color (4, 2, 1) (8, 0)
        8'b01101010, // Color (7, 3, 2) (9, 0)
        8'b00110110, // Color (3, 2, 1) (10, 0)
        8'b00111110, // Color (12, 9, 6) (11, 0)
        8'b00111110, // Color (12, 9, 6) (12, 0)
        8'b00111110, // Color (12, 9, 6) (13, 0)
        8'b00111010, // Color (11, 9, 5) (14, 0)
        8'b01101000, // Color (1, 1, 0) (15, 0)
        8'b01101000, // Color (1, 1, 0) (0, 1)
        8'b00111010, // Color (11, 9, 5) (1, 1)
        8'b00111100, // Color (10, 8, 5) (2, 1)
        8'b00111100, // Color (10, 8, 5) (3, 1)
        8'b00110100, // Color (9, 7, 4) (4, 1)
        8'b01000010, // Color (9, 8, 4) (5, 1)
        8'b00110110, // Color (3, 2, 1) (6, 1)
        8'b01011010, // Color (4, 2, 1) (7, 1)
        8'b01011010, // Color (4, 2, 1) (8, 1)
        8'b00110110, // Color (3, 2, 1) (9, 1)
        8'b00111100, // Color (10, 8, 5) (10, 1)
        8'b00111100, // Color (10, 8, 5) (11, 1)
        8'b00111010, // Color (11, 9, 5) (12, 1)
        8'b00111010, // Color (11, 9, 5) (13, 1)
        8'b01000010, // Color (9, 8, 4) (14, 1)
        8'b01101000, // Color (1, 1, 0) (15, 1)
        8'b01101000, // Color (1, 1, 0) (0, 2)
        8'b00111010, // Color (11, 9, 5) (1, 2)
        8'b00111010, // Color (11, 9, 5) (2, 2)
        8'b00111010, // Color (11, 9, 5) (3, 2)
        8'b00111100, // Color (10, 8, 5) (4, 2)
        8'b00111010, // Color (11, 9, 5) (5, 2)
        8'b00111100, // Color (10, 8, 5) (6, 2)
        8'b01110110, // Color (2, 2, 1) (7, 2)
        8'b01110110, // Color (2, 2, 1) (8, 2)
        8'b01000010, // Color (9, 8, 4) (9, 2)
        8'b01000010, // Color (9, 8, 4) (10, 2)
        8'b00111100, // Color (10, 8, 5) (11, 2)
        8'b00111100, // Color (10, 8, 5) (12, 2)
        8'b00111010, // Color (11, 9, 5) (13, 2)
        8'b00111010, // Color (11, 9, 5) (14, 2)
        8'b01101000, // Color (1, 1, 0) (15, 2)
        8'b01101000, // Color (1, 1, 0) (0, 3)
        8'b01000000, // Color (7, 6, 3) (1, 3)
        8'b01000000, // Color (7, 6, 3) (2, 3)
        8'b00110100, // Color (9, 7, 4) (3, 3)
        8'b00110100, // Color (9, 7, 4) (4, 3)
        8'b01000000, // Color (7, 6, 3) (5, 3)
        8'b01000100, // Color (6, 5, 2) (6, 3)
        8'b01101000, // Color (1, 1, 0) (7, 3)
        8'b01101000, // Color (1, 1, 0) (8, 3)
        8'b01000000, // Color (7, 6, 3) (9, 3)
        8'b01000100, // Color (6, 5, 2) (10, 3)
        8'b01000000, // Color (7, 6, 3) (11, 3)
        8'b01000100, // Color (6, 5, 2) (12, 3)
        8'b01000100, // Color (6, 5, 2) (13, 3)
        8'b01000000, // Color (7, 6, 3) (14, 3)
        8'b01101000, // Color (1, 1, 0) (15, 3)
        8'b01101000, // Color (1, 1, 0) (0, 4)
        8'b00111110, // Color (12, 9, 6) (1, 4)
        8'b01000010, // Color (9, 8, 4) (2, 4)
        8'b00111110, // Color (12, 9, 6) (3, 4)
        8'b00111110, // Color (12, 9, 6) (4, 4)
        8'b00111110, // Color (12, 9, 6) (5, 4)
        8'b00111110, // Color (12, 9, 6) (6, 4)
        8'b01011010, // Color (4, 2, 1) (7, 4)
        8'b01011010, // Color (4, 2, 1) (8, 4)
        8'b00111110, // Color (12, 9, 6) (9, 4)
        8'b00111110, // Color (12, 9, 6) (10, 4)
        8'b00111010, // Color (11, 9, 5) (11, 4)
        8'b00111100, // Color (10, 8, 5) (12, 4)
        8'b00111100, // Color (10, 8, 5) (13, 4)
        8'b01000010, // Color (9, 8, 4) (14, 4)
        8'b01101000, // Color (1, 1, 0) (15, 4)
        8'b01101000, // Color (1, 1, 0) (0, 5)
        8'b00111010, // Color (11, 9, 5) (1, 5)
        8'b00111010, // Color (11, 9, 5) (2, 5)
        8'b01101100, // Color (4, 2, 0) (3, 5)
        8'b01000010, // Color (9, 8, 4) (4, 5)
        8'b01101100, // Color (4, 2, 0) (5, 5)
        8'b01000010, // Color (9, 8, 4) (6, 5)
        8'b00110110, // Color (3, 2, 1) (7, 5)
        8'b00110110, // Color (3, 2, 1) (8, 5)
        8'b00111100, // Color (10, 8, 5) (9, 5)
        8'b00111100, // Color (10, 8, 5) (10, 5)
        8'b00111010, // Color (11, 9, 5) (11, 5)
        8'b00111010, // Color (11, 9, 5) (12, 5)
        8'b00111010, // Color (11, 9, 5) (13, 5)
        8'b00111010, // Color (11, 9, 5) (14, 5)
        8'b01101000, // Color (1, 1, 0) (15, 5)
        8'b01101000, // Color (1, 1, 0) (0, 6)
        8'b01000010, // Color (9, 8, 4) (1, 6)
        8'b00111100, // Color (10, 8, 5) (2, 6)
        8'b01101110, // Color (2, 1, 0) (3, 6)
        8'b00111100, // Color (10, 8, 5) (4, 6)
        8'b01101110, // Color (2, 1, 0) (5, 6)
        8'b00111100, // Color (10, 8, 5) (6, 6)
        8'b00110110, // Color (3, 2, 1) (7, 6)
        8'b00110110, // Color (3, 2, 1) (8, 6)
        8'b00111010, // Color (11, 9, 5) (9, 6)
        8'b00111010, // Color (11, 9, 5) (10, 6)
        8'b00111100, // Color (10, 8, 5) (11, 6)
        8'b00111100, // Color (10, 8, 5) (12, 6)
        8'b01000010, // Color (9, 8, 4) (13, 6)
        8'b01000010, // Color (9, 8, 4) (14, 6)
        8'b01101000, // Color (1, 1, 0) (15, 6)
        8'b01101000, // Color (1, 1, 0) (0, 7)
        8'b01000100, // Color (6, 5, 2) (1, 7)
        8'b01000000, // Color (7, 6, 3) (2, 7)
        8'b01000000, // Color (7, 6, 3) (3, 7)
        8'b01110010, // Color (13, 13, 13) (4, 7)
        8'b01000000, // Color (7, 6, 3) (5, 7)
        8'b01000100, // Color (6, 5, 2) (6, 7)
        8'b01101000, // Color (1, 1, 0) (7, 7)
        8'b01101000, // Color (1, 1, 0) (8, 7)
        8'b01000100, // Color (6, 5, 2) (9, 7)
        8'b01000000, // Color (7, 6, 3) (10, 7)
        8'b01000000, // Color (7, 6, 3) (11, 7)
        8'b01000000, // Color (7, 6, 3) (12, 7)
        8'b00110100, // Color (9, 7, 4) (13, 7)
        8'b01000000, // Color (7, 6, 3) (14, 7)
        8'b01101000, // Color (1, 1, 0) (15, 7)
        8'b01101000, // Color (1, 1, 0) (0, 8)
        8'b00111110, // Color (12, 9, 6) (1, 8)
        8'b00111110, // Color (12, 9, 6) (2, 8)
        8'b01110010, // Color (13, 13, 13) (3, 8)
        8'b00111100, // Color (10, 8, 5) (4, 8)
        8'b01110010, // Color (13, 13, 13) (5, 8)
        8'b00111110, // Color (12, 9, 6) (6, 8)
        8'b01011010, // Color (4, 2, 1) (7, 8)
        8'b01011010, // Color (4, 2, 1) (8, 8)
        8'b00111110, // Color (12, 9, 6) (9, 8)
        8'b00111110, // Color (12, 9, 6) (10, 8)
        8'b00111110, // Color (12, 9, 6) (11, 8)
        8'b00111110, // Color (12, 9, 6) (12, 8)
        8'b00111110, // Color (12, 9, 6) (13, 8)
        8'b00111010, // Color (11, 9, 5) (14, 8)
        8'b01101000, // Color (1, 1, 0) (15, 8)
        8'b01101000, // Color (1, 1, 0) (0, 9)
        8'b00111100, // Color (10, 8, 5) (1, 9)
        8'b00111010, // Color (11, 9, 5) (2, 9)
        8'b01100110, // Color (11, 11, 11) (3, 9)
        8'b00111010, // Color (11, 9, 5) (4, 9)
        8'b01100110, // Color (11, 11, 11) (5, 9)
        8'b00111100, // Color (10, 8, 5) (6, 9)
        8'b00110110, // Color (3, 2, 1) (7, 9)
        8'b00110110, // Color (3, 2, 1) (8, 9)
        8'b01000010, // Color (9, 8, 4) (9, 9)
        8'b00111100, // Color (10, 8, 5) (10, 9)
        8'b01000010, // Color (9, 8, 4) (11, 9)
        8'b00111100, // Color (10, 8, 5) (12, 9)
        8'b01000010, // Color (9, 8, 4) (13, 9)
        8'b01000010, // Color (9, 8, 4) (14, 9)
        8'b01101000, // Color (1, 1, 0) (15, 9)
        8'b01101000, // Color (1, 1, 0) (0, 10)
        8'b00111010, // Color (11, 9, 5) (1, 10)
        8'b00111100, // Color (10, 8, 5) (2, 10)
        8'b00111100, // Color (10, 8, 5) (3, 10)
        8'b01000010, // Color (9, 8, 4) (4, 10)
        8'b01000010, // Color (9, 8, 4) (5, 10)
        8'b01000010, // Color (9, 8, 4) (6, 10)
        8'b00110110, // Color (3, 2, 1) (7, 10)
        8'b00110110, // Color (3, 2, 1) (8, 10)
        8'b00111100, // Color (10, 8, 5) (9, 10)
        8'b00111100, // Color (10, 8, 5) (10, 10)
        8'b00111100, // Color (10, 8, 5) (11, 10)
        8'b01000010, // Color (9, 8, 4) (12, 10)
        8'b01000010, // Color (9, 8, 4) (13, 10)
        8'b00111010, // Color (11, 9, 5) (14, 10)
        8'b01101000, // Color (1, 1, 0) (15, 10)
        8'b01101000, // Color (1, 1, 0) (0, 11)
        8'b01000100, // Color (6, 5, 2) (1, 11)
        8'b01000000, // Color (7, 6, 3) (2, 11)
        8'b00110100, // Color (9, 7, 4) (3, 11)
        8'b00110100, // Color (9, 7, 4) (4, 11)
        8'b01000000, // Color (7, 6, 3) (5, 11)
        8'b01000100, // Color (6, 5, 2) (6, 11)
        8'b01110100, // Color (1, 0, 0) (7, 11)
        8'b01110100, // Color (1, 0, 0) (8, 11)
        8'b01000000, // Color (7, 6, 3) (9, 11)
        8'b00110100, // Color (9, 7, 4) (10, 11)
        8'b01000000, // Color (7, 6, 3) (11, 11)
        8'b01000000, // Color (7, 6, 3) (12, 11)
        8'b01000100, // Color (6, 5, 2) (13, 11)
        8'b01000100, // Color (6, 5, 2) (14, 11)
        8'b01101000, // Color (1, 1, 0) (15, 11)
        8'b01101000, // Color (1, 1, 0) (0, 12)
        8'b01000010, // Color (9, 8, 4) (1, 12)
        8'b00111010, // Color (11, 9, 5) (2, 12)
        8'b00111110, // Color (12, 9, 6) (3, 12)
        8'b00111110, // Color (12, 9, 6) (4, 12)
        8'b00111010, // Color (11, 9, 5) (5, 12)
        8'b00111010, // Color (11, 9, 5) (6, 12)
        8'b01011010, // Color (4, 2, 1) (7, 12)
        8'b01011010, // Color (4, 2, 1) (8, 12)
        8'b00111110, // Color (12, 9, 6) (9, 12)
        8'b00111110, // Color (12, 9, 6) (10, 12)
        8'b01000010, // Color (9, 8, 4) (11, 12)
        8'b00111110, // Color (12, 9, 6) (12, 12)
        8'b00111010, // Color (11, 9, 5) (13, 12)
        8'b00111110, // Color (12, 9, 6) (14, 12)
        8'b01101000, // Color (1, 1, 0) (15, 12)
        8'b01101000, // Color (1, 1, 0) (0, 13)
        8'b00111100, // Color (10, 8, 5) (1, 13)
        8'b00111010, // Color (11, 9, 5) (2, 13)
        8'b00111010, // Color (11, 9, 5) (3, 13)
        8'b01000010, // Color (9, 8, 4) (4, 13)
        8'b01000010, // Color (9, 8, 4) (5, 13)
        8'b00111100, // Color (10, 8, 5) (6, 13)
        8'b00110110, // Color (3, 2, 1) (7, 13)
        8'b00110110, // Color (3, 2, 1) (8, 13)
        8'b00111010, // Color (11, 9, 5) (9, 13)
        8'b00111010, // Color (11, 9, 5) (10, 13)
        8'b00111100, // Color (10, 8, 5) (11, 13)
        8'b00111010, // Color (11, 9, 5) (12, 13)
        8'b00111100, // Color (10, 8, 5) (13, 13)
        8'b00111100, // Color (10, 8, 5) (14, 13)
        8'b01101000, // Color (1, 1, 0) (15, 13)
        8'b01101000, // Color (1, 1, 0) (0, 14)
        8'b01000010, // Color (9, 8, 4) (1, 14)
        8'b01000010, // Color (9, 8, 4) (2, 14)
        8'b00111100, // Color (10, 8, 5) (3, 14)
        8'b00111010, // Color (11, 9, 5) (4, 14)
        8'b00111100, // Color (10, 8, 5) (5, 14)
        8'b01000010, // Color (9, 8, 4) (6, 14)
        8'b00110110, // Color (3, 2, 1) (7, 14)
        8'b00110110, // Color (3, 2, 1) (8, 14)
        8'b00111010, // Color (11, 9, 5) (9, 14)
        8'b00111100, // Color (10, 8, 5) (10, 14)
        8'b01000010, // Color (9, 8, 4) (11, 14)
        8'b01000010, // Color (9, 8, 4) (12, 14)
        8'b01000010, // Color (9, 8, 4) (13, 14)
        8'b01000010, // Color (9, 8, 4) (14, 14)
        8'b01101000, // Color (1, 1, 0) (15, 14)
        8'b01101000, // Color (1, 1, 0) (0, 15)
        8'b01000000, // Color (7, 6, 3) (1, 15)
        8'b01000000, // Color (7, 6, 3) (2, 15)
        8'b01000100, // Color (6, 5, 2) (3, 15)
        8'b01000100, // Color (6, 5, 2) (4, 15)
        8'b01000000, // Color (7, 6, 3) (5, 15)
        8'b00110100, // Color (9, 7, 4) (6, 15)
        8'b01101000, // Color (1, 1, 0) (7, 15)
        8'b01101000, // Color (1, 1, 0) (8, 15)
        8'b01000000, // Color (7, 6, 3) (9, 15)
        8'b01000100, // Color (6, 5, 2) (10, 15)
        8'b01000000, // Color (7, 6, 3) (11, 15)
        8'b01000100, // Color (6, 5, 2) (12, 15)
        8'b01000100, // Color (6, 5, 2) (13, 15)
        8'b01000100, // Color (6, 5, 2) (14, 15)
        8'b01101000, // Color (1, 1, 0) (15, 15)
        // 13_crafting_table_top
        8'b01101000, // Color (1, 1, 0) (0, 0)
        8'b01001000, // Color (0, 0, 0) (1, 0)
        8'b01001000, // Color (0, 0, 0) (2, 0)
        8'b01101000, // Color (1, 1, 0) (3, 0)
        8'b01101100, // Color (4, 2, 0) (4, 0)
        8'b01101010, // Color (7, 3, 2) (5, 0)
        8'b01101010, // Color (7, 3, 2) (6, 0)
        8'b01101010, // Color (7, 3, 2) (7, 0)
        8'b01101010, // Color (7, 3, 2) (8, 0)
        8'b01101010, // Color (7, 3, 2) (9, 0)
        8'b01101010, // Color (7, 3, 2) (10, 0)
        8'b01101100, // Color (4, 2, 0) (11, 0)
        8'b01101000, // Color (1, 1, 0) (12, 0)
        8'b01001000, // Color (0, 0, 0) (13, 0)
        8'b01101000, // Color (1, 1, 0) (14, 0)
        8'b01101000, // Color (1, 1, 0) (15, 0)
        8'b01001000, // Color (0, 0, 0) (0, 1)
        8'b01111000, // Color (11, 9, 6) (1, 1)
        8'b01111000, // Color (11, 9, 6) (2, 1)
        8'b01101100, // Color (4, 2, 0) (3, 1)
        8'b01111010, // Color (9, 5, 3) (4, 1)
        8'b01111100, // Color (10, 6, 3) (5, 1)
        8'b01111100, // Color (10, 6, 3) (6, 1)
        8'b01111100, // Color (10, 6, 3) (7, 1)
        8'b01111100, // Color (10, 6, 3) (8, 1)
        8'b01111100, // Color (10, 6, 3) (9, 1)
        8'b01111100, // Color (10, 6, 3) (10, 1)
        8'b01111010, // Color (9, 5, 3) (11, 1)
        8'b01101100, // Color (4, 2, 0) (12, 1)
        8'b01111000, // Color (11, 9, 6) (13, 1)
        8'b01111000, // Color (11, 9, 6) (14, 1)
        8'b01001000, // Color (0, 0, 0) (15, 1)
        8'b01001000, // Color (0, 0, 0) (0, 2)
        8'b01111000, // Color (11, 9, 6) (1, 2)
        8'b01101100, // Color (4, 2, 0) (2, 2)
        8'b01111100, // Color (10, 6, 3) (3, 2)
        8'b01111100, // Color (10, 6, 3) (4, 2)
        8'b01111100, // Color (10, 6, 3) (5, 2)
        8'b01111100, // Color (10, 6, 3) (6, 2)
        8'b01111100, // Color (10, 6, 3) (7, 2)
        8'b01111100, // Color (10, 6, 3) (8, 2)
        8'b01111100, // Color (10, 6, 3) (9, 2)
        8'b01111100, // Color (10, 6, 3) (10, 2)
        8'b01111100, // Color (10, 6, 3) (11, 2)
        8'b01111100, // Color (10, 6, 3) (12, 2)
        8'b01101100, // Color (4, 2, 0) (13, 2)
        8'b01111000, // Color (11, 9, 6) (14, 2)
        8'b01001000, // Color (0, 0, 0) (15, 2)
        8'b01101000, // Color (1, 1, 0) (0, 3)
        8'b01101100, // Color (4, 2, 0) (1, 3)
        8'b01111100, // Color (10, 6, 3) (2, 3)
        8'b00001000, // Color (5, 3, 2) (3, 3)
        8'b01011010, // Color (4, 2, 1) (4, 3)
        8'b00001000, // Color (5, 3, 2) (5, 3)
        8'b00001000, // Color (5, 3, 2) (6, 3)
        8'b00001000, // Color (5, 3, 2) (7, 3)
        8'b01011010, // Color (4, 2, 1) (8, 3)
        8'b01011010, // Color (4, 2, 1) (9, 3)
        8'b01011010, // Color (4, 2, 1) (10, 3)
        8'b01011010, // Color (4, 2, 1) (11, 3)
        8'b00001000, // Color (5, 3, 2) (12, 3)
        8'b01111100, // Color (10, 6, 3) (13, 3)
        8'b01101100, // Color (4, 2, 0) (14, 3)
        8'b01101000, // Color (1, 1, 0) (15, 3)
        8'b01101100, // Color (4, 2, 0) (0, 4)
        8'b01111010, // Color (9, 5, 3) (1, 4)
        8'b01111100, // Color (10, 6, 3) (2, 4)
        8'b00001000, // Color (5, 3, 2) (3, 4)
        8'b01111010, // Color (9, 5, 3) (4, 4)
        8'b01111100, // Color (10, 6, 3) (5, 4)
        8'b00001000, // Color (5, 3, 2) (6, 4)
        8'b01111100, // Color (10, 6, 3) (7, 4)
        8'b01111100, // Color (10, 6, 3) (8, 4)
        8'b01011010, // Color (4, 2, 1) (9, 4)
        8'b01111100, // Color (10, 6, 3) (10, 4)
        8'b01111100, // Color (10, 6, 3) (11, 4)
        8'b00001000, // Color (5, 3, 2) (12, 4)
        8'b01111100, // Color (10, 6, 3) (13, 4)
        8'b01111010, // Color (9, 5, 3) (14, 4)
        8'b01101100, // Color (4, 2, 0) (15, 4)
        8'b01101010, // Color (7, 3, 2) (0, 5)
        8'b01111100, // Color (10, 6, 3) (1, 5)
        8'b01111100, // Color (10, 6, 3) (2, 5)
        8'b00001000, // Color (5, 3, 2) (3, 5)
        8'b01111100, // Color (10, 6, 3) (4, 5)
        8'b01111100, // Color (10, 6, 3) (5, 5)
        8'b01011010, // Color (4, 2, 1) (6, 5)
        8'b01111010, // Color (9, 5, 3) (7, 5)
        8'b01111100, // Color (10, 6, 3) (8, 5)
        8'b00001000, // Color (5, 3, 2) (9, 5)
        8'b01111010, // Color (9, 5, 3) (10, 5)
        8'b01111100, // Color (10, 6, 3) (11, 5)
        8'b00001000, // Color (5, 3, 2) (12, 5)
        8'b01111100, // Color (10, 6, 3) (13, 5)
        8'b01111100, // Color (10, 6, 3) (14, 5)
        8'b01101010, // Color (7, 3, 2) (15, 5)
        8'b01101010, // Color (7, 3, 2) (0, 6)
        8'b01111100, // Color (10, 6, 3) (1, 6)
        8'b01111100, // Color (10, 6, 3) (2, 6)
        8'b00001000, // Color (5, 3, 2) (3, 6)
        8'b00001000, // Color (5, 3, 2) (4, 6)
        8'b01011010, // Color (4, 2, 1) (5, 6)
        8'b00001000, // Color (5, 3, 2) (6, 6)
        8'b00001000, // Color (5, 3, 2) (7, 6)
        8'b01011010, // Color (4, 2, 1) (8, 6)
        8'b00001000, // Color (5, 3, 2) (9, 6)
        8'b00001000, // Color (5, 3, 2) (10, 6)
        8'b01011010, // Color (4, 2, 1) (11, 6)
        8'b00001000, // Color (5, 3, 2) (12, 6)
        8'b01111100, // Color (10, 6, 3) (13, 6)
        8'b01111100, // Color (10, 6, 3) (14, 6)
        8'b01101010, // Color (7, 3, 2) (15, 6)
        8'b01101010, // Color (7, 3, 2) (0, 7)
        8'b01111100, // Color (10, 6, 3) (1, 7)
        8'b01111100, // Color (10, 6, 3) (2, 7)
        8'b00001000, // Color (5, 3, 2) (3, 7)
        8'b01111100, // Color (10, 6, 3) (4, 7)
        8'b01111100, // Color (10, 6, 3) (5, 7)
        8'b00001000, // Color (5, 3, 2) (6, 7)
        8'b01111100, // Color (10, 6, 3) (7, 7)
        8'b01111100, // Color (10, 6, 3) (8, 7)
        8'b00001000, // Color (5, 3, 2) (9, 7)
        8'b01111100, // Color (10, 6, 3) (10, 7)
        8'b01111100, // Color (10, 6, 3) (11, 7)
        8'b00001000, // Color (5, 3, 2) (12, 7)
        8'b01111100, // Color (10, 6, 3) (13, 7)
        8'b01111100, // Color (10, 6, 3) (14, 7)
        8'b01101010, // Color (7, 3, 2) (15, 7)
        8'b01101010, // Color (7, 3, 2) (0, 8)
        8'b01111100, // Color (10, 6, 3) (1, 8)
        8'b01111100, // Color (10, 6, 3) (2, 8)
        8'b00001000, // Color (5, 3, 2) (3, 8)
        8'b01111100, // Color (10, 6, 3) (4, 8)
        8'b01111100, // Color (10, 6, 3) (5, 8)
        8'b00001000, // Color (5, 3, 2) (6, 8)
        8'b01111100, // Color (10, 6, 3) (7, 8)
        8'b01111100, // Color (10, 6, 3) (8, 8)
        8'b00001000, // Color (5, 3, 2) (9, 8)
        8'b01111100, // Color (10, 6, 3) (10, 8)
        8'b01111100, // Color (10, 6, 3) (11, 8)
        8'b00001000, // Color (5, 3, 2) (12, 8)
        8'b01111100, // Color (10, 6, 3) (13, 8)
        8'b01111100, // Color (10, 6, 3) (14, 8)
        8'b01101010, // Color (7, 3, 2) (15, 8)
        8'b01101010, // Color (7, 3, 2) (0, 9)
        8'b01111100, // Color (10, 6, 3) (1, 9)
        8'b01111100, // Color (10, 6, 3) (2, 9)
        8'b01011010, // Color (4, 2, 1) (3, 9)
        8'b01011010, // Color (4, 2, 1) (4, 9)
        8'b01011010, // Color (4, 2, 1) (5, 9)
        8'b00001000, // Color (5, 3, 2) (6, 9)
        8'b01011010, // Color (4, 2, 1) (7, 9)
        8'b01011010, // Color (4, 2, 1) (8, 9)
        8'b00001000, // Color (5, 3, 2) (9, 9)
        8'b00001000, // Color (5, 3, 2) (10, 9)
        8'b01011010, // Color (4, 2, 1) (11, 9)
        8'b00001000, // Color (5, 3, 2) (12, 9)
        8'b01111100, // Color (10, 6, 3) (13, 9)
        8'b01111100, // Color (10, 6, 3) (14, 9)
        8'b01101010, // Color (7, 3, 2) (15, 9)
        8'b01101010, // Color (7, 3, 2) (0, 10)
        8'b01111100, // Color (10, 6, 3) (1, 10)
        8'b01111100, // Color (10, 6, 3) (2, 10)
        8'b01011010, // Color (4, 2, 1) (3, 10)
        8'b01111010, // Color (9, 5, 3) (4, 10)
        8'b01111100, // Color (10, 6, 3) (5, 10)
        8'b01011010, // Color (4, 2, 1) (6, 10)
        8'b01111100, // Color (10, 6, 3) (7, 10)
        8'b01111010, // Color (9, 5, 3) (8, 10)
        8'b01011010, // Color (4, 2, 1) (9, 10)
        8'b01111100, // Color (10, 6, 3) (10, 10)
        8'b01111100, // Color (10, 6, 3) (11, 10)
        8'b00001000, // Color (5, 3, 2) (12, 10)
        8'b01111100, // Color (10, 6, 3) (13, 10)
        8'b01111100, // Color (10, 6, 3) (14, 10)
        8'b01101010, // Color (7, 3, 2) (15, 10)
        8'b01101100, // Color (4, 2, 0) (0, 11)
        8'b01111010, // Color (9, 5, 3) (1, 11)
        8'b01111100, // Color (10, 6, 3) (2, 11)
        8'b00001000, // Color (5, 3, 2) (3, 11)
        8'b01111010, // Color (9, 5, 3) (4, 11)
        8'b01111100, // Color (10, 6, 3) (5, 11)
        8'b01011010, // Color (4, 2, 1) (6, 11)
        8'b01111100, // Color (10, 6, 3) (7, 11)
        8'b01111100, // Color (10, 6, 3) (8, 11)
        8'b01011010, // Color (4, 2, 1) (9, 11)
        8'b01111010, // Color (9, 5, 3) (10, 11)
        8'b01111100, // Color (10, 6, 3) (11, 11)
        8'b00001000, // Color (5, 3, 2) (12, 11)
        8'b01111100, // Color (10, 6, 3) (13, 11)
        8'b01111010, // Color (9, 5, 3) (14, 11)
        8'b01101100, // Color (4, 2, 0) (15, 11)
        8'b01101000, // Color (1, 1, 0) (0, 12)
        8'b01101100, // Color (4, 2, 0) (1, 12)
        8'b01111100, // Color (10, 6, 3) (2, 12)
        8'b00001000, // Color (5, 3, 2) (3, 12)
        8'b00001000, // Color (5, 3, 2) (4, 12)
        8'b01011010, // Color (4, 2, 1) (5, 12)
        8'b00001000, // Color (5, 3, 2) (6, 12)
        8'b00001000, // Color (5, 3, 2) (7, 12)
        8'b00001000, // Color (5, 3, 2) (8, 12)
        8'b00001000, // Color (5, 3, 2) (9, 12)
        8'b00001000, // Color (5, 3, 2) (10, 12)
        8'b00001000, // Color (5, 3, 2) (11, 12)
        8'b00001000, // Color (5, 3, 2) (12, 12)
        8'b01111100, // Color (10, 6, 3) (13, 12)
        8'b01101100, // Color (4, 2, 0) (14, 12)
        8'b01101000, // Color (1, 1, 0) (15, 12)
        8'b01001000, // Color (0, 0, 0) (0, 13)
        8'b01111000, // Color (11, 9, 6) (1, 13)
        8'b01101100, // Color (4, 2, 0) (2, 13)
        8'b01111100, // Color (10, 6, 3) (3, 13)
        8'b01111100, // Color (10, 6, 3) (4, 13)
        8'b01111100, // Color (10, 6, 3) (5, 13)
        8'b01111100, // Color (10, 6, 3) (6, 13)
        8'b01111100, // Color (10, 6, 3) (7, 13)
        8'b01111100, // Color (10, 6, 3) (8, 13)
        8'b01111100, // Color (10, 6, 3) (9, 13)
        8'b01111100, // Color (10, 6, 3) (10, 13)
        8'b01111100, // Color (10, 6, 3) (11, 13)
        8'b01111100, // Color (10, 6, 3) (12, 13)
        8'b01101100, // Color (4, 2, 0) (13, 13)
        8'b01111000, // Color (11, 9, 6) (14, 13)
        8'b01001000, // Color (0, 0, 0) (15, 13)
        8'b01101000, // Color (1, 1, 0) (0, 14)
        8'b01111000, // Color (11, 9, 6) (1, 14)
        8'b01111000, // Color (11, 9, 6) (2, 14)
        8'b01101100, // Color (4, 2, 0) (3, 14)
        8'b01111010, // Color (9, 5, 3) (4, 14)
        8'b01111100, // Color (10, 6, 3) (5, 14)
        8'b01111100, // Color (10, 6, 3) (6, 14)
        8'b01111100, // Color (10, 6, 3) (7, 14)
        8'b01111100, // Color (10, 6, 3) (8, 14)
        8'b01111100, // Color (10, 6, 3) (9, 14)
        8'b01111100, // Color (10, 6, 3) (10, 14)
        8'b01111010, // Color (9, 5, 3) (11, 14)
        8'b01101100, // Color (4, 2, 0) (12, 14)
        8'b01111000, // Color (11, 9, 6) (13, 14)
        8'b01111000, // Color (11, 9, 6) (14, 14)
        8'b01101000, // Color (1, 1, 0) (15, 14)
        8'b01101000, // Color (1, 1, 0) (0, 15)
        8'b01101000, // Color (1, 1, 0) (1, 15)
        8'b01001000, // Color (0, 0, 0) (2, 15)
        8'b01101000, // Color (1, 1, 0) (3, 15)
        8'b01101100, // Color (4, 2, 0) (4, 15)
        8'b01101010, // Color (7, 3, 2) (5, 15)
        8'b01101010, // Color (7, 3, 2) (6, 15)
        8'b01101010, // Color (7, 3, 2) (7, 15)
        8'b01101010, // Color (7, 3, 2) (8, 15)
        8'b01101010, // Color (7, 3, 2) (9, 15)
        8'b01101010, // Color (7, 3, 2) (10, 15)
        8'b01101100, // Color (4, 2, 0) (11, 15)
        8'b01101000, // Color (1, 1, 0) (12, 15)
        8'b01001000, // Color (0, 0, 0) (13, 15)
        8'b01001000, // Color (0, 0, 0) (14, 15)
        8'b01101000, // Color (1, 1, 0) (15, 15)
        // 14_iron_block
        8'b01111110, // Color (13, 12, 12) (0, 0)
        8'b10000000, // Color (12, 12, 12) (1, 0)
        8'b10000000, // Color (12, 12, 12) (2, 0)
        8'b01111110, // Color (13, 12, 12) (3, 0)
        8'b01111110, // Color (13, 12, 12) (4, 0)
        8'b01111110, // Color (13, 12, 12) (5, 0)
        8'b01111110, // Color (13, 12, 12) (6, 0)
        8'b01111110, // Color (13, 12, 12) (7, 0)
        8'b01111110, // Color (13, 12, 12) (8, 0)
        8'b01111110, // Color (13, 12, 12) (9, 0)
        8'b01111110, // Color (13, 12, 12) (10, 0)
        8'b10000000, // Color (12, 12, 12) (11, 0)
        8'b10000000, // Color (12, 12, 12) (12, 0)
        8'b10000000, // Color (12, 12, 12) (13, 0)
        8'b10000000, // Color (12, 12, 12) (14, 0)
        8'b01111110, // Color (13, 12, 12) (15, 0)
        8'b10000000, // Color (12, 12, 12) (0, 1)
        8'b01110000, // Color (15, 15, 15) (1, 1)
        8'b01110000, // Color (15, 15, 15) (2, 1)
        8'b01110000, // Color (15, 15, 15) (3, 1)
        8'b01110000, // Color (15, 15, 15) (4, 1)
        8'b01110000, // Color (15, 15, 15) (5, 1)
        8'b10000010, // Color (14, 14, 14) (6, 1)
        8'b10000010, // Color (14, 14, 14) (7, 1)
        8'b10000010, // Color (14, 14, 14) (8, 1)
        8'b10000010, // Color (14, 14, 14) (9, 1)
        8'b10000010, // Color (14, 14, 14) (10, 1)
        8'b10000010, // Color (14, 14, 14) (11, 1)
        8'b10000010, // Color (14, 14, 14) (12, 1)
        8'b10000010, // Color (14, 14, 14) (13, 1)
        8'b10000010, // Color (14, 14, 14) (14, 1)
        8'b10000000, // Color (12, 12, 12) (15, 1)
        8'b10000000, // Color (12, 12, 12) (0, 2)
        8'b10000010, // Color (14, 14, 14) (1, 2)
        8'b10000010, // Color (14, 14, 14) (2, 2)
        8'b10000010, // Color (14, 14, 14) (3, 2)
        8'b10000010, // Color (14, 14, 14) (4, 2)
        8'b10000010, // Color (14, 14, 14) (5, 2)
        8'b10000010, // Color (14, 14, 14) (6, 2)
        8'b10000010, // Color (14, 14, 14) (7, 2)
        8'b10000010, // Color (14, 14, 14) (8, 2)
        8'b10000010, // Color (14, 14, 14) (9, 2)
        8'b10000010, // Color (14, 14, 14) (10, 2)
        8'b10000010, // Color (14, 14, 14) (11, 2)
        8'b10000010, // Color (14, 14, 14) (12, 2)
        8'b10000010, // Color (14, 14, 14) (13, 2)
        8'b10000010, // Color (14, 14, 14) (14, 2)
        8'b01100110, // Color (11, 11, 11) (15, 2)
        8'b01100110, // Color (11, 11, 11) (0, 3)
        8'b01110010, // Color (13, 13, 13) (1, 3)
        8'b01110010, // Color (13, 13, 13) (2, 3)
        8'b01110010, // Color (13, 13, 13) (3, 3)
        8'b01110010, // Color (13, 13, 13) (4, 3)
        8'b01110010, // Color (13, 13, 13) (5, 3)
        8'b01110010, // Color (13, 13, 13) (6, 3)
        8'b01110010, // Color (13, 13, 13) (7, 3)
        8'b10000010, // Color (14, 14, 14) (8, 3)
        8'b10000010, // Color (14, 14, 14) (9, 3)
        8'b10000010, // Color (14, 14, 14) (10, 3)
        8'b01110010, // Color (13, 13, 13) (11, 3)
        8'b01110010, // Color (13, 13, 13) (12, 3)
        8'b01110010, // Color (13, 13, 13) (13, 3)
        8'b01110010, // Color (13, 13, 13) (14, 3)
        8'b01100110, // Color (11, 11, 11) (15, 3)
        8'b10000000, // Color (12, 12, 12) (0, 4)
        8'b01110000, // Color (15, 15, 15) (1, 4)
        8'b01110000, // Color (15, 15, 15) (2, 4)
        8'b01110000, // Color (15, 15, 15) (3, 4)
        8'b01110000, // Color (15, 15, 15) (4, 4)
        8'b01110000, // Color (15, 15, 15) (5, 4)
        8'b01110000, // Color (15, 15, 15) (6, 4)
        8'b10000010, // Color (14, 14, 14) (7, 4)
        8'b10000010, // Color (14, 14, 14) (8, 4)
        8'b10000010, // Color (14, 14, 14) (9, 4)
        8'b10000010, // Color (14, 14, 14) (10, 4)
        8'b10000010, // Color (14, 14, 14) (11, 4)
        8'b10000010, // Color (14, 14, 14) (12, 4)
        8'b10000010, // Color (14, 14, 14) (13, 4)
        8'b10000010, // Color (14, 14, 14) (14, 4)
        8'b01100110, // Color (11, 11, 11) (15, 4)
        8'b10000000, // Color (12, 12, 12) (0, 5)
        8'b10000010, // Color (14, 14, 14) (1, 5)
        8'b10000010, // Color (14, 14, 14) (2, 5)
        8'b10000010, // Color (14, 14, 14) (3, 5)
        8'b10000010, // Color (14, 14, 14) (4, 5)
        8'b10000010, // Color (14, 14, 14) (5, 5)
        8'b10000010, // Color (14, 14, 14) (6, 5)
        8'b10000010, // Color (14, 14, 14) (7, 5)
        8'b10000010, // Color (14, 14, 14) (8, 5)
        8'b10000010, // Color (14, 14, 14) (9, 5)
        8'b10000010, // Color (14, 14, 14) (10, 5)
        8'b10000010, // Color (14, 14, 14) (11, 5)
        8'b10000010, // Color (14, 14, 14) (12, 5)
        8'b10000010, // Color (14, 14, 14) (13, 5)
        8'b10000010, // Color (14, 14, 14) (14, 5)
        8'b01100110, // Color (11, 11, 11) (15, 5)
        8'b01100110, // Color (11, 11, 11) (0, 6)
        8'b01110010, // Color (13, 13, 13) (1, 6)
        8'b01110010, // Color (13, 13, 13) (2, 6)
        8'b01110010, // Color (13, 13, 13) (3, 6)
        8'b01110010, // Color (13, 13, 13) (4, 6)
        8'b01110010, // Color (13, 13, 13) (5, 6)
        8'b10000010, // Color (14, 14, 14) (6, 6)
        8'b10000010, // Color (14, 14, 14) (7, 6)
        8'b10000010, // Color (14, 14, 14) (8, 6)
        8'b10000010, // Color (14, 14, 14) (9, 6)
        8'b01110010, // Color (13, 13, 13) (10, 6)
        8'b01110010, // Color (13, 13, 13) (11, 6)
        8'b01110010, // Color (13, 13, 13) (12, 6)
        8'b01110010, // Color (13, 13, 13) (13, 6)
        8'b01110010, // Color (13, 13, 13) (14, 6)
        8'b01100110, // Color (11, 11, 11) (15, 6)
        8'b10000000, // Color (12, 12, 12) (0, 7)
        8'b01110000, // Color (15, 15, 15) (1, 7)
        8'b01110000, // Color (15, 15, 15) (2, 7)
        8'b10000010, // Color (14, 14, 14) (3, 7)
        8'b10000010, // Color (14, 14, 14) (4, 7)
        8'b10000010, // Color (14, 14, 14) (5, 7)
        8'b10000010, // Color (14, 14, 14) (6, 7)
        8'b10000010, // Color (14, 14, 14) (7, 7)
        8'b10000010, // Color (14, 14, 14) (8, 7)
        8'b10000010, // Color (14, 14, 14) (9, 7)
        8'b10000010, // Color (14, 14, 14) (10, 7)
        8'b10000010, // Color (14, 14, 14) (11, 7)
        8'b10000010, // Color (14, 14, 14) (12, 7)
        8'b10000010, // Color (14, 14, 14) (13, 7)
        8'b10000010, // Color (14, 14, 14) (14, 7)
        8'b01100110, // Color (11, 11, 11) (15, 7)
        8'b10000000, // Color (12, 12, 12) (0, 8)
        8'b10000010, // Color (14, 14, 14) (1, 8)
        8'b10000010, // Color (14, 14, 14) (2, 8)
        8'b10000010, // Color (14, 14, 14) (3, 8)
        8'b10000010, // Color (14, 14, 14) (4, 8)
        8'b10000010, // Color (14, 14, 14) (5, 8)
        8'b10000010, // Color (14, 14, 14) (6, 8)
        8'b10000010, // Color (14, 14, 14) (7, 8)
        8'b10000010, // Color (14, 14, 14) (8, 8)
        8'b10000010, // Color (14, 14, 14) (9, 8)
        8'b10000010, // Color (14, 14, 14) (10, 8)
        8'b10000010, // Color (14, 14, 14) (11, 8)
        8'b10000010, // Color (14, 14, 14) (12, 8)
        8'b10000010, // Color (14, 14, 14) (13, 8)
        8'b10000010, // Color (14, 14, 14) (14, 8)
        8'b01100110, // Color (11, 11, 11) (15, 8)
        8'b01100110, // Color (11, 11, 11) (0, 9)
        8'b01110010, // Color (13, 13, 13) (1, 9)
        8'b01110010, // Color (13, 13, 13) (2, 9)
        8'b01110010, // Color (13, 13, 13) (3, 9)
        8'b01110010, // Color (13, 13, 13) (4, 9)
        8'b01110010, // Color (13, 13, 13) (5, 9)
        8'b01110010, // Color (13, 13, 13) (6, 9)
        8'b01110010, // Color (13, 13, 13) (7, 9)
        8'b01110010, // Color (13, 13, 13) (8, 9)
        8'b10000010, // Color (14, 14, 14) (9, 9)
        8'b10000010, // Color (14, 14, 14) (10, 9)
        8'b10000010, // Color (14, 14, 14) (11, 9)
        8'b01110010, // Color (13, 13, 13) (12, 9)
        8'b01110010, // Color (13, 13, 13) (13, 9)
        8'b01110010, // Color (13, 13, 13) (14, 9)
        8'b01100110, // Color (11, 11, 11) (15, 9)
        8'b10000000, // Color (12, 12, 12) (0, 10)
        8'b01110000, // Color (15, 15, 15) (1, 10)
        8'b01110000, // Color (15, 15, 15) (2, 10)
        8'b01110000, // Color (15, 15, 15) (3, 10)
        8'b01110000, // Color (15, 15, 15) (4, 10)
        8'b01110000, // Color (15, 15, 15) (5, 10)
        8'b01110000, // Color (15, 15, 15) (6, 10)
        8'b10000010, // Color (14, 14, 14) (7, 10)
        8'b10000010, // Color (14, 14, 14) (8, 10)
        8'b10000010, // Color (14, 14, 14) (9, 10)
        8'b10000010, // Color (14, 14, 14) (10, 10)
        8'b10000010, // Color (14, 14, 14) (11, 10)
        8'b10000010, // Color (14, 14, 14) (12, 10)
        8'b10000010, // Color (14, 14, 14) (13, 10)
        8'b10000010, // Color (14, 14, 14) (14, 10)
        8'b01100110, // Color (11, 11, 11) (15, 10)
        8'b10000000, // Color (12, 12, 12) (0, 11)
        8'b10000010, // Color (14, 14, 14) (1, 11)
        8'b10000010, // Color (14, 14, 14) (2, 11)
        8'b10000010, // Color (14, 14, 14) (3, 11)
        8'b10000010, // Color (14, 14, 14) (4, 11)
        8'b10000010, // Color (14, 14, 14) (5, 11)
        8'b10000010, // Color (14, 14, 14) (6, 11)
        8'b10000010, // Color (14, 14, 14) (7, 11)
        8'b10000010, // Color (14, 14, 14) (8, 11)
        8'b10000010, // Color (14, 14, 14) (9, 11)
        8'b10000010, // Color (14, 14, 14) (10, 11)
        8'b10000010, // Color (14, 14, 14) (11, 11)
        8'b10000010, // Color (14, 14, 14) (12, 11)
        8'b10000010, // Color (14, 14, 14) (13, 11)
        8'b10000010, // Color (14, 14, 14) (14, 11)
        8'b01100110, // Color (11, 11, 11) (15, 11)
        8'b01100110, // Color (11, 11, 11) (0, 12)
        8'b01110010, // Color (13, 13, 13) (1, 12)
        8'b01110010, // Color (13, 13, 13) (2, 12)
        8'b01110010, // Color (13, 13, 13) (3, 12)
        8'b01110010, // Color (13, 13, 13) (4, 12)
        8'b01110010, // Color (13, 13, 13) (5, 12)
        8'b01110010, // Color (13, 13, 13) (6, 12)
        8'b10000010, // Color (14, 14, 14) (7, 12)
        8'b10000010, // Color (14, 14, 14) (8, 12)
        8'b10000010, // Color (14, 14, 14) (9, 12)
        8'b10000010, // Color (14, 14, 14) (10, 12)
        8'b01110010, // Color (13, 13, 13) (11, 12)
        8'b01110010, // Color (13, 13, 13) (12, 12)
        8'b01110010, // Color (13, 13, 13) (13, 12)
        8'b01110010, // Color (13, 13, 13) (14, 12)
        8'b01100110, // Color (11, 11, 11) (15, 12)
        8'b10000000, // Color (12, 12, 12) (0, 13)
        8'b01110000, // Color (15, 15, 15) (1, 13)
        8'b01110000, // Color (15, 15, 15) (2, 13)
        8'b01110000, // Color (15, 15, 15) (3, 13)
        8'b01110000, // Color (15, 15, 15) (4, 13)
        8'b10000010, // Color (14, 14, 14) (5, 13)
        8'b10000010, // Color (14, 14, 14) (6, 13)
        8'b10000010, // Color (14, 14, 14) (7, 13)
        8'b10000010, // Color (14, 14, 14) (8, 13)
        8'b10000010, // Color (14, 14, 14) (9, 13)
        8'b10000010, // Color (14, 14, 14) (10, 13)
        8'b10000010, // Color (14, 14, 14) (11, 13)
        8'b10000010, // Color (14, 14, 14) (12, 13)
        8'b10000010, // Color (14, 14, 14) (13, 13)
        8'b10000010, // Color (14, 14, 14) (14, 13)
        8'b01100110, // Color (11, 11, 11) (15, 13)
        8'b10000000, // Color (12, 12, 12) (0, 14)
        8'b10000010, // Color (14, 14, 14) (1, 14)
        8'b10000010, // Color (14, 14, 14) (2, 14)
        8'b10000010, // Color (14, 14, 14) (3, 14)
        8'b10000010, // Color (14, 14, 14) (4, 14)
        8'b10000010, // Color (14, 14, 14) (5, 14)
        8'b10000010, // Color (14, 14, 14) (6, 14)
        8'b10000010, // Color (14, 14, 14) (7, 14)
        8'b10000010, // Color (14, 14, 14) (8, 14)
        8'b10000010, // Color (14, 14, 14) (9, 14)
        8'b10000010, // Color (14, 14, 14) (10, 14)
        8'b10000010, // Color (14, 14, 14) (11, 14)
        8'b10000010, // Color (14, 14, 14) (12, 14)
        8'b10000010, // Color (14, 14, 14) (13, 14)
        8'b10000010, // Color (14, 14, 14) (14, 14)
        8'b01100110, // Color (11, 11, 11) (15, 14)
        8'b10000000, // Color (12, 12, 12) (0, 15)
        8'b10000000, // Color (12, 12, 12) (1, 15)
        8'b10000000, // Color (12, 12, 12) (2, 15)
        8'b10000000, // Color (12, 12, 12) (3, 15)
        8'b10000000, // Color (12, 12, 12) (4, 15)
        8'b10000000, // Color (12, 12, 12) (5, 15)
        8'b10000000, // Color (12, 12, 12) (6, 15)
        8'b01100110, // Color (11, 11, 11) (7, 15)
        8'b01100110, // Color (11, 11, 11) (8, 15)
        8'b10000000, // Color (12, 12, 12) (9, 15)
        8'b01100110, // Color (11, 11, 11) (10, 15)
        8'b01100110, // Color (11, 11, 11) (11, 15)
        8'b01100110, // Color (11, 11, 11) (12, 15)
        8'b01100110, // Color (11, 11, 11) (13, 15)
        8'b01100110, // Color (11, 11, 11) (14, 15)
        8'b01100110, // Color (11, 11, 11) (15, 15)
        // 15_gold_block
        8'b10000100, // Color (15, 12, 2) (0, 0)
        8'b10000100, // Color (15, 12, 2) (1, 0)
        8'b10000100, // Color (15, 12, 2) (2, 0)
        8'b10000100, // Color (15, 12, 2) (3, 0)
        8'b10000110, // Color (15, 11, 2) (4, 0)
        8'b10000110, // Color (15, 11, 2) (5, 0)
        8'b10000100, // Color (15, 12, 2) (6, 0)
        8'b10000100, // Color (15, 12, 2) (7, 0)
        8'b10000100, // Color (15, 12, 2) (8, 0)
        8'b10000110, // Color (15, 11, 2) (9, 0)
        8'b10000110, // Color (15, 11, 2) (10, 0)
        8'b10000110, // Color (15, 11, 2) (11, 0)
        8'b10000110, // Color (15, 11, 2) (12, 0)
        8'b10000100, // Color (15, 12, 2) (13, 0)
        8'b10000100, // Color (15, 12, 2) (14, 0)
        8'b10001000, // Color (13, 9, 3) (15, 0)
        8'b10000100, // Color (15, 12, 2) (0, 1)
        8'b10001010, // Color (15, 15, 9) (1, 1)
        8'b10001100, // Color (15, 15, 11) (2, 1)
        8'b10001100, // Color (15, 15, 11) (3, 1)
        8'b10001110, // Color (15, 14, 4) (4, 1)
        8'b10001110, // Color (15, 14, 4) (5, 1)
        8'b10001010, // Color (15, 15, 9) (6, 1)
        8'b10001010, // Color (15, 15, 9) (7, 1)
        8'b10001010, // Color (15, 15, 9) (8, 1)
        8'b10001110, // Color (15, 14, 4) (9, 1)
        8'b10001110, // Color (15, 14, 4) (10, 1)
        8'b10010000, // Color (15, 13, 3) (11, 1)
        8'b10010000, // Color (15, 13, 3) (12, 1)
        8'b10001010, // Color (15, 15, 9) (13, 1)
        8'b10001010, // Color (15, 15, 9) (14, 1)
        8'b10001000, // Color (13, 9, 3) (15, 1)
        8'b10000100, // Color (15, 12, 2) (0, 2)
        8'b10001100, // Color (15, 15, 11) (1, 2)
        8'b10010000, // Color (15, 13, 3) (2, 2)
        8'b10010000, // Color (15, 13, 3) (3, 2)
        8'b10001110, // Color (15, 14, 4) (4, 2)
        8'b10001010, // Color (15, 15, 9) (5, 2)
        8'b10001110, // Color (15, 14, 4) (6, 2)
        8'b10001110, // Color (15, 14, 4) (7, 2)
        8'b10010000, // Color (15, 13, 3) (8, 2)
        8'b10000100, // Color (15, 12, 2) (9, 2)
        8'b10000110, // Color (15, 11, 2) (10, 2)
        8'b10000110, // Color (15, 11, 2) (11, 2)
        8'b10000100, // Color (15, 12, 2) (12, 2)
        8'b10001110, // Color (15, 14, 4) (13, 2)
        8'b10001010, // Color (15, 15, 9) (14, 2)
        8'b10001000, // Color (13, 9, 3) (15, 2)
        8'b10000100, // Color (15, 12, 2) (0, 3)
        8'b10001100, // Color (15, 15, 11) (1, 3)
        8'b10010000, // Color (15, 13, 3) (2, 3)
        8'b10001110, // Color (15, 14, 4) (3, 3)
        8'b10001010, // Color (15, 15, 9) (4, 3)
        8'b10001110, // Color (15, 14, 4) (5, 3)
        8'b10001110, // Color (15, 14, 4) (6, 3)
        8'b10001110, // Color (15, 14, 4) (7, 3)
        8'b10010000, // Color (15, 13, 3) (8, 3)
        8'b10000100, // Color (15, 12, 2) (9, 3)
        8'b10000100, // Color (15, 12, 2) (10, 3)
        8'b10000100, // Color (15, 12, 2) (11, 3)
        8'b10001110, // Color (15, 14, 4) (12, 3)
        8'b10001110, // Color (15, 14, 4) (13, 3)
        8'b10001110, // Color (15, 14, 4) (14, 3)
        8'b10001000, // Color (13, 9, 3) (15, 3)
        8'b10000110, // Color (15, 11, 2) (0, 4)
        8'b10001110, // Color (15, 14, 4) (1, 4)
        8'b10001110, // Color (15, 14, 4) (2, 4)
        8'b10001110, // Color (15, 14, 4) (3, 4)
        8'b10001110, // Color (15, 14, 4) (4, 4)
        8'b10001110, // Color (15, 14, 4) (5, 4)
        8'b10001110, // Color (15, 14, 4) (6, 4)
        8'b10010000, // Color (15, 13, 3) (7, 4)
        8'b10000100, // Color (15, 12, 2) (8, 4)
        8'b10000100, // Color (15, 12, 2) (9, 4)
        8'b10010000, // Color (15, 13, 3) (10, 4)
        8'b10001110, // Color (15, 14, 4) (11, 4)
        8'b10001110, // Color (15, 14, 4) (12, 4)
        8'b10010000, // Color (15, 13, 3) (13, 4)
        8'b10001110, // Color (15, 14, 4) (14, 4)
        8'b10001000, // Color (13, 9, 3) (15, 4)
        8'b10000110, // Color (15, 11, 2) (0, 5)
        8'b10001110, // Color (15, 14, 4) (1, 5)
        8'b10001110, // Color (15, 14, 4) (2, 5)
        8'b10001110, // Color (15, 14, 4) (3, 5)
        8'b10001110, // Color (15, 14, 4) (4, 5)
        8'b10001110, // Color (15, 14, 4) (5, 5)
        8'b10010000, // Color (15, 13, 3) (6, 5)
        8'b10000100, // Color (15, 12, 2) (7, 5)
        8'b10000100, // Color (15, 12, 2) (8, 5)
        8'b10010000, // Color (15, 13, 3) (9, 5)
        8'b10001110, // Color (15, 14, 4) (10, 5)
        8'b10001110, // Color (15, 14, 4) (11, 5)
        8'b10010000, // Color (15, 13, 3) (12, 5)
        8'b10000100, // Color (15, 12, 2) (13, 5)
        8'b10000110, // Color (15, 11, 2) (14, 5)
        8'b10010010, // Color (12, 8, 2) (15, 5)
        8'b10000100, // Color (15, 12, 2) (0, 6)
        8'b10001010, // Color (15, 15, 9) (1, 6)
        8'b10001110, // Color (15, 14, 4) (2, 6)
        8'b10001110, // Color (15, 14, 4) (3, 6)
        8'b10001110, // Color (15, 14, 4) (4, 6)
        8'b10001110, // Color (15, 14, 4) (5, 6)
        8'b10001110, // Color (15, 14, 4) (6, 6)
        8'b10010000, // Color (15, 13, 3) (7, 6)
        8'b10010000, // Color (15, 13, 3) (8, 6)
        8'b10001110, // Color (15, 14, 4) (9, 6)
        8'b10001110, // Color (15, 14, 4) (10, 6)
        8'b10010000, // Color (15, 13, 3) (11, 6)
        8'b10000100, // Color (15, 12, 2) (12, 6)
        8'b10000110, // Color (15, 11, 2) (13, 6)
        8'b10000110, // Color (15, 11, 2) (14, 6)
        8'b10010010, // Color (12, 8, 2) (15, 6)
        8'b10000100, // Color (15, 12, 2) (0, 7)
        8'b10001010, // Color (15, 15, 9) (1, 7)
        8'b10001110, // Color (15, 14, 4) (2, 7)
        8'b10001110, // Color (15, 14, 4) (3, 7)
        8'b10001110, // Color (15, 14, 4) (4, 7)
        8'b10001110, // Color (15, 14, 4) (5, 7)
        8'b10010000, // Color (15, 13, 3) (6, 7)
        8'b10010000, // Color (15, 13, 3) (7, 7)
        8'b10001110, // Color (15, 14, 4) (8, 7)
        8'b10001110, // Color (15, 14, 4) (9, 7)
        8'b10010000, // Color (15, 13, 3) (10, 7)
        8'b10000100, // Color (15, 12, 2) (11, 7)
        8'b10000100, // Color (15, 12, 2) (12, 7)
        8'b10000110, // Color (15, 11, 2) (13, 7)
        8'b10000100, // Color (15, 12, 2) (14, 7)
        8'b10010010, // Color (12, 8, 2) (15, 7)
        8'b10000110, // Color (15, 11, 2) (0, 8)
        8'b10001110, // Color (15, 14, 4) (1, 8)
        8'b10001110, // Color (15, 14, 4) (2, 8)
        8'b10001110, // Color (15, 14, 4) (3, 8)
        8'b10001110, // Color (15, 14, 4) (4, 8)
        8'b10010000, // Color (15, 13, 3) (5, 8)
        8'b10010000, // Color (15, 13, 3) (6, 8)
        8'b10001110, // Color (15, 14, 4) (7, 8)
        8'b10001110, // Color (15, 14, 4) (8, 8)
        8'b10010000, // Color (15, 13, 3) (9, 8)
        8'b10010000, // Color (15, 13, 3) (10, 8)
        8'b10000100, // Color (15, 12, 2) (11, 8)
        8'b10000100, // Color (15, 12, 2) (12, 8)
        8'b10000100, // Color (15, 12, 2) (13, 8)
        8'b10010000, // Color (15, 13, 3) (14, 8)
        8'b10001000, // Color (13, 9, 3) (15, 8)
        8'b10000110, // Color (15, 11, 2) (0, 9)
        8'b10001110, // Color (15, 14, 4) (1, 9)
        8'b10001110, // Color (15, 14, 4) (2, 9)
        8'b10001110, // Color (15, 14, 4) (3, 9)
        8'b10010000, // Color (15, 13, 3) (4, 9)
        8'b10010000, // Color (15, 13, 3) (5, 9)
        8'b10001110, // Color (15, 14, 4) (6, 9)
        8'b10001110, // Color (15, 14, 4) (7, 9)
        8'b10010000, // Color (15, 13, 3) (8, 9)
        8'b10010000, // Color (15, 13, 3) (9, 9)
        8'b10010000, // Color (15, 13, 3) (10, 9)
        8'b10010000, // Color (15, 13, 3) (11, 9)
        8'b10000100, // Color (15, 12, 2) (12, 9)
        8'b10001110, // Color (15, 14, 4) (13, 9)
        8'b10010000, // Color (15, 13, 3) (14, 9)
        8'b10001000, // Color (13, 9, 3) (15, 9)
        8'b10000110, // Color (15, 11, 2) (0, 10)
        8'b10010000, // Color (15, 13, 3) (1, 10)
        8'b10001110, // Color (15, 14, 4) (2, 10)
        8'b10010000, // Color (15, 13, 3) (3, 10)
        8'b10010000, // Color (15, 13, 3) (4, 10)
        8'b10001110, // Color (15, 14, 4) (5, 10)
        8'b10001110, // Color (15, 14, 4) (6, 10)
        8'b10010000, // Color (15, 13, 3) (7, 10)
        8'b10010000, // Color (15, 13, 3) (8, 10)
        8'b10010000, // Color (15, 13, 3) (9, 10)
        8'b10010000, // Color (15, 13, 3) (10, 10)
        8'b10010000, // Color (15, 13, 3) (11, 10)
        8'b10001110, // Color (15, 14, 4) (12, 10)
        8'b10001110, // Color (15, 14, 4) (13, 10)
        8'b10000100, // Color (15, 12, 2) (14, 10)
        8'b10010010, // Color (12, 8, 2) (15, 10)
        8'b10000110, // Color (15, 11, 2) (0, 11)
        8'b10000100, // Color (15, 12, 2) (1, 11)
        8'b10010000, // Color (15, 13, 3) (2, 11)
        8'b10010000, // Color (15, 13, 3) (3, 11)
        8'b10001110, // Color (15, 14, 4) (4, 11)
        8'b10001110, // Color (15, 14, 4) (5, 11)
        8'b10010000, // Color (15, 13, 3) (6, 11)
        8'b10000100, // Color (15, 12, 2) (7, 11)
        8'b10000100, // Color (15, 12, 2) (8, 11)
        8'b10010000, // Color (15, 13, 3) (9, 11)
        8'b10000100, // Color (15, 12, 2) (10, 11)
        8'b10001110, // Color (15, 14, 4) (11, 11)
        8'b10001110, // Color (15, 14, 4) (12, 11)
        8'b10010000, // Color (15, 13, 3) (13, 11)
        8'b10000100, // Color (15, 12, 2) (14, 11)
        8'b10010010, // Color (12, 8, 2) (15, 11)
        8'b10000110, // Color (15, 11, 2) (0, 12)
        8'b10000100, // Color (15, 12, 2) (1, 12)
        8'b10010000, // Color (15, 13, 3) (2, 12)
        8'b10001110, // Color (15, 14, 4) (3, 12)
        8'b10001110, // Color (15, 14, 4) (4, 12)
        8'b10010000, // Color (15, 13, 3) (5, 12)
        8'b10000100, // Color (15, 12, 2) (6, 12)
        8'b10000110, // Color (15, 11, 2) (7, 12)
        8'b10000110, // Color (15, 11, 2) (8, 12)
        8'b10000100, // Color (15, 12, 2) (9, 12)
        8'b10001110, // Color (15, 14, 4) (10, 12)
        8'b10001110, // Color (15, 14, 4) (11, 12)
        8'b10010000, // Color (15, 13, 3) (12, 12)
        8'b10000100, // Color (15, 12, 2) (13, 12)
        8'b10010000, // Color (15, 13, 3) (14, 12)
        8'b10001000, // Color (13, 9, 3) (15, 12)
        8'b10000110, // Color (15, 11, 2) (0, 13)
        8'b10000110, // Color (15, 11, 2) (1, 13)
        8'b10001110, // Color (15, 14, 4) (2, 13)
        8'b10001110, // Color (15, 14, 4) (3, 13)
        8'b10010000, // Color (15, 13, 3) (4, 13)
        8'b10000100, // Color (15, 12, 2) (5, 13)
        8'b10000110, // Color (15, 11, 2) (6, 13)
        8'b10000110, // Color (15, 11, 2) (7, 13)
        8'b10000100, // Color (15, 12, 2) (8, 13)
        8'b10010000, // Color (15, 13, 3) (9, 13)
        8'b10010000, // Color (15, 13, 3) (10, 13)
        8'b10010000, // Color (15, 13, 3) (11, 13)
        8'b10000100, // Color (15, 12, 2) (12, 13)
        8'b10000100, // Color (15, 12, 2) (13, 13)
        8'b10001110, // Color (15, 14, 4) (14, 13)
        8'b10001000, // Color (13, 9, 3) (15, 13)
        8'b10000110, // Color (15, 11, 2) (0, 14)
        8'b10000100, // Color (15, 12, 2) (1, 14)
        8'b10000110, // Color (15, 11, 2) (2, 14)
        8'b10000100, // Color (15, 12, 2) (3, 14)
        8'b10000100, // Color (15, 12, 2) (4, 14)
        8'b10000110, // Color (15, 11, 2) (5, 14)
        8'b10000110, // Color (15, 11, 2) (6, 14)
        8'b10000100, // Color (15, 12, 2) (7, 14)
        8'b10010000, // Color (15, 13, 3) (8, 14)
        8'b10010000, // Color (15, 13, 3) (9, 14)
        8'b10000100, // Color (15, 12, 2) (10, 14)
        8'b10000100, // Color (15, 12, 2) (11, 14)
        8'b10010000, // Color (15, 13, 3) (12, 14)
        8'b10001110, // Color (15, 14, 4) (13, 14)
        8'b10001110, // Color (15, 14, 4) (14, 14)
        8'b10010010, // Color (12, 8, 2) (15, 14)
        8'b10001000, // Color (13, 9, 3) (0, 15)
        8'b10001000, // Color (13, 9, 3) (1, 15)
        8'b10010010, // Color (12, 8, 2) (2, 15)
        8'b10001000, // Color (13, 9, 3) (3, 15)
        8'b10001000, // Color (13, 9, 3) (4, 15)
        8'b10010010, // Color (12, 8, 2) (5, 15)
        8'b10010010, // Color (12, 8, 2) (6, 15)
        8'b10010010, // Color (12, 8, 2) (7, 15)
        8'b10001000, // Color (13, 9, 3) (8, 15)
        8'b10001000, // Color (13, 9, 3) (9, 15)
        8'b10010010, // Color (12, 8, 2) (10, 15)
        8'b10010010, // Color (12, 8, 2) (11, 15)
        8'b10001000, // Color (13, 9, 3) (12, 15)
        8'b10001000, // Color (13, 9, 3) (13, 15)
        8'b10010010, // Color (12, 8, 2) (14, 15)
        8'b10010010, // Color (12, 8, 2) (15, 15)
        // 16_redstone_block
        8'b10010100, // Color (14, 2, 0) (0, 0)
        8'b10010100, // Color (14, 2, 0) (1, 0)
        8'b10010100, // Color (14, 2, 0) (2, 0)
        8'b10010100, // Color (14, 2, 0) (3, 0)
        8'b10010100, // Color (14, 2, 0) (4, 0)
        8'b10010100, // Color (14, 2, 0) (5, 0)
        8'b10010100, // Color (14, 2, 0) (6, 0)
        8'b10010100, // Color (14, 2, 0) (7, 0)
        8'b10010100, // Color (14, 2, 0) (8, 0)
        8'b10010100, // Color (14, 2, 0) (9, 0)
        8'b10010100, // Color (14, 2, 0) (10, 0)
        8'b10010100, // Color (14, 2, 0) (11, 0)
        8'b10010100, // Color (14, 2, 0) (12, 0)
        8'b10010100, // Color (14, 2, 0) (13, 0)
        8'b10010100, // Color (14, 2, 0) (14, 0)
        8'b10010100, // Color (14, 2, 0) (15, 0)
        8'b10010100, // Color (14, 2, 0) (0, 1)
        8'b10010110, // Color (11, 2, 0) (1, 1)
        8'b10010110, // Color (11, 2, 0) (2, 1)
        8'b10010100, // Color (14, 2, 0) (3, 1)
        8'b10010110, // Color (11, 2, 0) (4, 1)
        8'b10010110, // Color (11, 2, 0) (5, 1)
        8'b10011000, // Color (10, 1, 0) (6, 1)
        8'b10011000, // Color (10, 1, 0) (7, 1)
        8'b10011000, // Color (10, 1, 0) (8, 1)
        8'b10010110, // Color (11, 2, 0) (9, 1)
        8'b10010110, // Color (11, 2, 0) (10, 1)
        8'b10010100, // Color (14, 2, 0) (11, 1)
        8'b10010110, // Color (11, 2, 0) (12, 1)
        8'b10010110, // Color (11, 2, 0) (13, 1)
        8'b10010110, // Color (11, 2, 0) (14, 1)
        8'b10010100, // Color (14, 2, 0) (15, 1)
        8'b10010100, // Color (14, 2, 0) (0, 2)
        8'b10010110, // Color (11, 2, 0) (1, 2)
        8'b10010110, // Color (11, 2, 0) (2, 2)
        8'b10010100, // Color (14, 2, 0) (3, 2)
        8'b10011000, // Color (10, 1, 0) (4, 2)
        8'b10011000, // Color (10, 1, 0) (5, 2)
        8'b10011010, // Color (7, 0, 0) (6, 2)
        8'b10011000, // Color (10, 1, 0) (7, 2)
        8'b10011000, // Color (10, 1, 0) (8, 2)
        8'b10011000, // Color (10, 1, 0) (9, 2)
        8'b10011000, // Color (10, 1, 0) (10, 2)
        8'b10011000, // Color (10, 1, 0) (11, 2)
        8'b10010110, // Color (11, 2, 0) (12, 2)
        8'b10011000, // Color (10, 1, 0) (13, 2)
        8'b10010110, // Color (11, 2, 0) (14, 2)
        8'b10010100, // Color (14, 2, 0) (15, 2)
        8'b10010100, // Color (14, 2, 0) (0, 3)
        8'b10010110, // Color (11, 2, 0) (1, 3)
        8'b10010110, // Color (11, 2, 0) (2, 3)
        8'b10011000, // Color (10, 1, 0) (3, 3)
        8'b10010110, // Color (11, 2, 0) (4, 3)
        8'b10011100, // Color (9, 1, 0) (5, 3)
        8'b10011100, // Color (9, 1, 0) (6, 3)
        8'b10011010, // Color (7, 0, 0) (7, 3)
        8'b10011010, // Color (7, 0, 0) (8, 3)
        8'b10011100, // Color (9, 1, 0) (9, 3)
        8'b10011100, // Color (9, 1, 0) (10, 3)
        8'b10011000, // Color (10, 1, 0) (11, 3)
        8'b10011010, // Color (7, 0, 0) (12, 3)
        8'b10011000, // Color (10, 1, 0) (13, 3)
        8'b10010110, // Color (11, 2, 0) (14, 3)
        8'b10010100, // Color (14, 2, 0) (15, 3)
        8'b10010100, // Color (14, 2, 0) (0, 4)
        8'b10010100, // Color (14, 2, 0) (1, 4)
        8'b10010110, // Color (11, 2, 0) (2, 4)
        8'b10011000, // Color (10, 1, 0) (3, 4)
        8'b10011100, // Color (9, 1, 0) (4, 4)
        8'b10011100, // Color (9, 1, 0) (5, 4)
        8'b10011010, // Color (7, 0, 0) (6, 4)
        8'b10011100, // Color (9, 1, 0) (7, 4)
        8'b10011000, // Color (10, 1, 0) (8, 4)
        8'b10011010, // Color (7, 0, 0) (9, 4)
        8'b10011100, // Color (9, 1, 0) (10, 4)
        8'b10011100, // Color (9, 1, 0) (11, 4)
        8'b10011000, // Color (10, 1, 0) (12, 4)
        8'b10010100, // Color (14, 2, 0) (13, 4)
        8'b10010100, // Color (14, 2, 0) (14, 4)
        8'b10010100, // Color (14, 2, 0) (15, 4)
        8'b10010100, // Color (14, 2, 0) (0, 5)
        8'b10010110, // Color (11, 2, 0) (1, 5)
        8'b10011000, // Color (10, 1, 0) (2, 5)
        8'b10011100, // Color (9, 1, 0) (3, 5)
        8'b10011010, // Color (7, 0, 0) (4, 5)
        8'b10011010, // Color (7, 0, 0) (5, 5)
        8'b10011010, // Color (7, 0, 0) (6, 5)
        8'b10011010, // Color (7, 0, 0) (7, 5)
        8'b10011010, // Color (7, 0, 0) (8, 5)
        8'b10011010, // Color (7, 0, 0) (9, 5)
        8'b10011010, // Color (7, 0, 0) (10, 5)
        8'b10011010, // Color (7, 0, 0) (11, 5)
        8'b10010100, // Color (14, 2, 0) (12, 5)
        8'b10011000, // Color (10, 1, 0) (13, 5)
        8'b10010110, // Color (11, 2, 0) (14, 5)
        8'b10010100, // Color (14, 2, 0) (15, 5)
        8'b10010100, // Color (14, 2, 0) (0, 6)
        8'b10010110, // Color (11, 2, 0) (1, 6)
        8'b10011010, // Color (7, 0, 0) (2, 6)
        8'b10011000, // Color (10, 1, 0) (3, 6)
        8'b10011100, // Color (9, 1, 0) (4, 6)
        8'b10011010, // Color (7, 0, 0) (5, 6)
        8'b10011010, // Color (7, 0, 0) (6, 6)
        8'b10011010, // Color (7, 0, 0) (7, 6)
        8'b10011010, // Color (7, 0, 0) (8, 6)
        8'b10011010, // Color (7, 0, 0) (9, 6)
        8'b10011010, // Color (7, 0, 0) (10, 6)
        8'b10011100, // Color (9, 1, 0) (11, 6)
        8'b10011100, // Color (9, 1, 0) (12, 6)
        8'b10011100, // Color (9, 1, 0) (13, 6)
        8'b10010110, // Color (11, 2, 0) (14, 6)
        8'b10010100, // Color (14, 2, 0) (15, 6)
        8'b10010100, // Color (14, 2, 0) (0, 7)
        8'b10011000, // Color (10, 1, 0) (1, 7)
        8'b10011100, // Color (9, 1, 0) (2, 7)
        8'b10011100, // Color (9, 1, 0) (3, 7)
        8'b10011010, // Color (7, 0, 0) (4, 7)
        8'b10011010, // Color (7, 0, 0) (5, 7)
        8'b10011010, // Color (7, 0, 0) (6, 7)
        8'b10011010, // Color (7, 0, 0) (7, 7)
        8'b10011010, // Color (7, 0, 0) (8, 7)
        8'b10011010, // Color (7, 0, 0) (9, 7)
        8'b10011010, // Color (7, 0, 0) (10, 7)
        8'b10011010, // Color (7, 0, 0) (11, 7)
        8'b10011100, // Color (9, 1, 0) (12, 7)
        8'b10011000, // Color (10, 1, 0) (13, 7)
        8'b10011000, // Color (10, 1, 0) (14, 7)
        8'b10010100, // Color (14, 2, 0) (15, 7)
        8'b10010100, // Color (14, 2, 0) (0, 8)
        8'b10011000, // Color (10, 1, 0) (1, 8)
        8'b10011000, // Color (10, 1, 0) (2, 8)
        8'b10010110, // Color (11, 2, 0) (3, 8)
        8'b10011100, // Color (9, 1, 0) (4, 8)
        8'b10011010, // Color (7, 0, 0) (5, 8)
        8'b10011010, // Color (7, 0, 0) (6, 8)
        8'b10011010, // Color (7, 0, 0) (7, 8)
        8'b10011010, // Color (7, 0, 0) (8, 8)
        8'b10011010, // Color (7, 0, 0) (9, 8)
        8'b10011010, // Color (7, 0, 0) (10, 8)
        8'b10011100, // Color (9, 1, 0) (11, 8)
        8'b10011100, // Color (9, 1, 0) (12, 8)
        8'b10011100, // Color (9, 1, 0) (13, 8)
        8'b10010110, // Color (11, 2, 0) (14, 8)
        8'b10010100, // Color (14, 2, 0) (15, 8)
        8'b10010100, // Color (14, 2, 0) (0, 9)
        8'b10010110, // Color (11, 2, 0) (1, 9)
        8'b10011000, // Color (10, 1, 0) (2, 9)
        8'b10010100, // Color (14, 2, 0) (3, 9)
        8'b10011100, // Color (9, 1, 0) (4, 9)
        8'b10011100, // Color (9, 1, 0) (5, 9)
        8'b10011010, // Color (7, 0, 0) (6, 9)
        8'b10011000, // Color (10, 1, 0) (7, 9)
        8'b10011100, // Color (9, 1, 0) (8, 9)
        8'b10011010, // Color (7, 0, 0) (9, 9)
        8'b10011100, // Color (9, 1, 0) (10, 9)
        8'b10011100, // Color (9, 1, 0) (11, 9)
        8'b10011100, // Color (9, 1, 0) (12, 9)
        8'b10011000, // Color (10, 1, 0) (13, 9)
        8'b10010110, // Color (11, 2, 0) (14, 9)
        8'b10010100, // Color (14, 2, 0) (15, 9)
        8'b10010100, // Color (14, 2, 0) (0, 10)
        8'b10010110, // Color (11, 2, 0) (1, 10)
        8'b10011000, // Color (10, 1, 0) (2, 10)
        8'b10011100, // Color (9, 1, 0) (3, 10)
        8'b10011100, // Color (9, 1, 0) (4, 10)
        8'b10011010, // Color (7, 0, 0) (5, 10)
        8'b10011010, // Color (7, 0, 0) (6, 10)
        8'b10011010, // Color (7, 0, 0) (7, 10)
        8'b10010100, // Color (14, 2, 0) (8, 10)
        8'b10011010, // Color (7, 0, 0) (9, 10)
        8'b10011010, // Color (7, 0, 0) (10, 10)
        8'b10011100, // Color (9, 1, 0) (11, 10)
        8'b10011000, // Color (10, 1, 0) (12, 10)
        8'b10011000, // Color (10, 1, 0) (13, 10)
        8'b10010100, // Color (14, 2, 0) (14, 10)
        8'b10010100, // Color (14, 2, 0) (15, 10)
        8'b10010100, // Color (14, 2, 0) (0, 11)
        8'b10010110, // Color (11, 2, 0) (1, 11)
        8'b10010110, // Color (11, 2, 0) (2, 11)
        8'b10011000, // Color (10, 1, 0) (3, 11)
        8'b10011100, // Color (9, 1, 0) (4, 11)
        8'b10011100, // Color (9, 1, 0) (5, 11)
        8'b10011010, // Color (7, 0, 0) (6, 11)
        8'b10011100, // Color (9, 1, 0) (7, 11)
        8'b10011010, // Color (7, 0, 0) (8, 11)
        8'b10011010, // Color (7, 0, 0) (9, 11)
        8'b10011100, // Color (9, 1, 0) (10, 11)
        8'b10011100, // Color (9, 1, 0) (11, 11)
        8'b10011100, // Color (9, 1, 0) (12, 11)
        8'b10011010, // Color (7, 0, 0) (13, 11)
        8'b10010110, // Color (11, 2, 0) (14, 11)
        8'b10010100, // Color (14, 2, 0) (15, 11)
        8'b10010100, // Color (14, 2, 0) (0, 12)
        8'b10010110, // Color (11, 2, 0) (1, 12)
        8'b10011000, // Color (10, 1, 0) (2, 12)
        8'b10011000, // Color (10, 1, 0) (3, 12)
        8'b10011000, // Color (10, 1, 0) (4, 12)
        8'b10011100, // Color (9, 1, 0) (5, 12)
        8'b10011100, // Color (9, 1, 0) (6, 12)
        8'b10011100, // Color (9, 1, 0) (7, 12)
        8'b10011100, // Color (9, 1, 0) (8, 12)
        8'b10011100, // Color (9, 1, 0) (9, 12)
        8'b10011100, // Color (9, 1, 0) (10, 12)
        8'b10011000, // Color (10, 1, 0) (11, 12)
        8'b10011000, // Color (10, 1, 0) (12, 12)
        8'b10011000, // Color (10, 1, 0) (13, 12)
        8'b10011000, // Color (10, 1, 0) (14, 12)
        8'b10010100, // Color (14, 2, 0) (15, 12)
        8'b10010100, // Color (14, 2, 0) (0, 13)
        8'b10010100, // Color (14, 2, 0) (1, 13)
        8'b10010110, // Color (11, 2, 0) (2, 13)
        8'b10011100, // Color (9, 1, 0) (3, 13)
        8'b10011000, // Color (10, 1, 0) (4, 13)
        8'b10010100, // Color (14, 2, 0) (5, 13)
        8'b10011000, // Color (10, 1, 0) (6, 13)
        8'b10011100, // Color (9, 1, 0) (7, 13)
        8'b10011100, // Color (9, 1, 0) (8, 13)
        8'b10011010, // Color (7, 0, 0) (9, 13)
        8'b10011000, // Color (10, 1, 0) (10, 13)
        8'b10011000, // Color (10, 1, 0) (11, 13)
        8'b10010110, // Color (11, 2, 0) (12, 13)
        8'b10011000, // Color (10, 1, 0) (13, 13)
        8'b10010110, // Color (11, 2, 0) (14, 13)
        8'b10010100, // Color (14, 2, 0) (15, 13)
        8'b10010100, // Color (14, 2, 0) (0, 14)
        8'b10010110, // Color (11, 2, 0) (1, 14)
        8'b10010110, // Color (11, 2, 0) (2, 14)
        8'b10010110, // Color (11, 2, 0) (3, 14)
        8'b10010100, // Color (14, 2, 0) (4, 14)
        8'b10010100, // Color (14, 2, 0) (5, 14)
        8'b10010110, // Color (11, 2, 0) (6, 14)
        8'b10010110, // Color (11, 2, 0) (7, 14)
        8'b10011000, // Color (10, 1, 0) (8, 14)
        8'b10011000, // Color (10, 1, 0) (9, 14)
        8'b10010110, // Color (11, 2, 0) (10, 14)
        8'b10010110, // Color (11, 2, 0) (11, 14)
        8'b10010110, // Color (11, 2, 0) (12, 14)
        8'b10010110, // Color (11, 2, 0) (13, 14)
        8'b10010110, // Color (11, 2, 0) (14, 14)
        8'b10010100, // Color (14, 2, 0) (15, 14)
        8'b10010100, // Color (14, 2, 0) (0, 15)
        8'b10010100, // Color (14, 2, 0) (1, 15)
        8'b10010100, // Color (14, 2, 0) (2, 15)
        8'b10010100, // Color (14, 2, 0) (3, 15)
        8'b10010100, // Color (14, 2, 0) (4, 15)
        8'b10010100, // Color (14, 2, 0) (5, 15)
        8'b10010100, // Color (14, 2, 0) (6, 15)
        8'b10010100, // Color (14, 2, 0) (7, 15)
        8'b10010100, // Color (14, 2, 0) (8, 15)
        8'b10010100, // Color (14, 2, 0) (9, 15)
        8'b10010100, // Color (14, 2, 0) (10, 15)
        8'b10010100, // Color (14, 2, 0) (11, 15)
        8'b10010100, // Color (14, 2, 0) (12, 15)
        8'b10010100, // Color (14, 2, 0) (13, 15)
        8'b10010100, // Color (14, 2, 0) (14, 15)
        8'b10010100, // Color (14, 2, 0) (15, 15)
        // 17_diamond_block
        8'b10011110, // Color (4, 14, 14) (0, 0)
        8'b10011110, // Color (4, 14, 14) (1, 0)
        8'b10011110, // Color (4, 14, 14) (2, 0)
        8'b10011110, // Color (4, 14, 14) (3, 0)
        8'b10100000, // Color (3, 14, 14) (4, 0)
        8'b10100000, // Color (3, 14, 14) (5, 0)
        8'b10011110, // Color (4, 14, 14) (6, 0)
        8'b10011110, // Color (4, 14, 14) (7, 0)
        8'b10011110, // Color (4, 14, 14) (8, 0)
        8'b10100000, // Color (3, 14, 14) (9, 0)
        8'b10100000, // Color (3, 14, 14) (10, 0)
        8'b10100000, // Color (3, 14, 14) (11, 0)
        8'b10100000, // Color (3, 14, 14) (12, 0)
        8'b10011110, // Color (4, 14, 14) (13, 0)
        8'b10011110, // Color (4, 14, 14) (14, 0)
        8'b10100010, // Color (1, 12, 12) (15, 0)
        8'b10011110, // Color (4, 14, 14) (0, 1)
        8'b10100100, // Color (13, 15, 15) (1, 1)
        8'b01110000, // Color (15, 15, 15) (2, 1)
        8'b01110000, // Color (15, 15, 15) (3, 1)
        8'b10100110, // Color (9, 15, 14) (4, 1)
        8'b10100110, // Color (9, 15, 14) (5, 1)
        8'b10100100, // Color (13, 15, 15) (6, 1)
        8'b10100100, // Color (13, 15, 15) (7, 1)
        8'b10100100, // Color (13, 15, 15) (8, 1)
        8'b10100110, // Color (9, 15, 14) (9, 1)
        8'b10100110, // Color (9, 15, 14) (10, 1)
        8'b10101000, // Color (6, 15, 14) (11, 1)
        8'b10101000, // Color (6, 15, 14) (12, 1)
        8'b10100100, // Color (13, 15, 15) (13, 1)
        8'b10100100, // Color (13, 15, 15) (14, 1)
        8'b10100010, // Color (1, 12, 12) (15, 1)
        8'b10011110, // Color (4, 14, 14) (0, 2)
        8'b01110000, // Color (15, 15, 15) (1, 2)
        8'b10101000, // Color (6, 15, 14) (2, 2)
        8'b10101000, // Color (6, 15, 14) (3, 2)
        8'b10101010, // Color (7, 15, 15) (4, 2)
        8'b10100100, // Color (13, 15, 15) (5, 2)
        8'b10100110, // Color (9, 15, 14) (6, 2)
        8'b10100110, // Color (9, 15, 14) (7, 2)
        8'b10101000, // Color (6, 15, 14) (8, 2)
        8'b10011110, // Color (4, 14, 14) (9, 2)
        8'b10100000, // Color (3, 14, 14) (10, 2)
        8'b10100000, // Color (3, 14, 14) (11, 2)
        8'b10011110, // Color (4, 14, 14) (12, 2)
        8'b10101010, // Color (7, 15, 15) (13, 2)
        8'b10100100, // Color (13, 15, 15) (14, 2)
        8'b10100010, // Color (1, 12, 12) (15, 2)
        8'b10011110, // Color (4, 14, 14) (0, 3)
        8'b01110000, // Color (15, 15, 15) (1, 3)
        8'b10101000, // Color (6, 15, 14) (2, 3)
        8'b10101010, // Color (7, 15, 15) (3, 3)
        8'b10100100, // Color (13, 15, 15) (4, 3)
        8'b10100110, // Color (9, 15, 14) (5, 3)
        8'b10100110, // Color (9, 15, 14) (6, 3)
        8'b10101010, // Color (7, 15, 15) (7, 3)
        8'b10101000, // Color (6, 15, 14) (8, 3)
        8'b10011110, // Color (4, 14, 14) (9, 3)
        8'b10011110, // Color (4, 14, 14) (10, 3)
        8'b10011110, // Color (4, 14, 14) (11, 3)
        8'b10101010, // Color (7, 15, 15) (12, 3)
        8'b10101010, // Color (7, 15, 15) (13, 3)
        8'b10100110, // Color (9, 15, 14) (14, 3)
        8'b10100010, // Color (1, 12, 12) (15, 3)
        8'b10100000, // Color (3, 14, 14) (0, 4)
        8'b10100110, // Color (9, 15, 14) (1, 4)
        8'b10101010, // Color (7, 15, 15) (2, 4)
        8'b10100110, // Color (9, 15, 14) (3, 4)
        8'b10100110, // Color (9, 15, 14) (4, 4)
        8'b10100110, // Color (9, 15, 14) (5, 4)
        8'b10101010, // Color (7, 15, 15) (6, 4)
        8'b10101000, // Color (6, 15, 14) (7, 4)
        8'b10011110, // Color (4, 14, 14) (8, 4)
        8'b10011110, // Color (4, 14, 14) (9, 4)
        8'b10101000, // Color (6, 15, 14) (10, 4)
        8'b10101010, // Color (7, 15, 15) (11, 4)
        8'b10101010, // Color (7, 15, 15) (12, 4)
        8'b10101000, // Color (6, 15, 14) (13, 4)
        8'b10100110, // Color (9, 15, 14) (14, 4)
        8'b10100010, // Color (1, 12, 12) (15, 4)
        8'b10100000, // Color (3, 14, 14) (0, 5)
        8'b10100110, // Color (9, 15, 14) (1, 5)
        8'b10100110, // Color (9, 15, 14) (2, 5)
        8'b10100110, // Color (9, 15, 14) (3, 5)
        8'b10100110, // Color (9, 15, 14) (4, 5)
        8'b10101010, // Color (7, 15, 15) (5, 5)
        8'b10101000, // Color (6, 15, 14) (6, 5)
        8'b10011110, // Color (4, 14, 14) (7, 5)
        8'b10011110, // Color (4, 14, 14) (8, 5)
        8'b10101000, // Color (6, 15, 14) (9, 5)
        8'b10100110, // Color (9, 15, 14) (10, 5)
        8'b10100110, // Color (9, 15, 14) (11, 5)
        8'b10101000, // Color (6, 15, 14) (12, 5)
        8'b10011110, // Color (4, 14, 14) (13, 5)
        8'b10100000, // Color (3, 14, 14) (14, 5)
        8'b10101100, // Color (0, 11, 11) (15, 5)
        8'b10011110, // Color (4, 14, 14) (0, 6)
        8'b10100100, // Color (13, 15, 15) (1, 6)
        8'b10100110, // Color (9, 15, 14) (2, 6)
        8'b10100110, // Color (9, 15, 14) (3, 6)
        8'b10101010, // Color (7, 15, 15) (4, 6)
        8'b10101010, // Color (7, 15, 15) (5, 6)
        8'b10101010, // Color (7, 15, 15) (6, 6)
        8'b10101000, // Color (6, 15, 14) (7, 6)
        8'b10101000, // Color (6, 15, 14) (8, 6)
        8'b10100110, // Color (9, 15, 14) (9, 6)
        8'b10100110, // Color (9, 15, 14) (10, 6)
        8'b10101000, // Color (6, 15, 14) (11, 6)
        8'b10011110, // Color (4, 14, 14) (12, 6)
        8'b10100000, // Color (3, 14, 14) (13, 6)
        8'b10100000, // Color (3, 14, 14) (14, 6)
        8'b10101100, // Color (0, 11, 11) (15, 6)
        8'b10011110, // Color (4, 14, 14) (0, 7)
        8'b10100100, // Color (13, 15, 15) (1, 7)
        8'b10100110, // Color (9, 15, 14) (2, 7)
        8'b10101010, // Color (7, 15, 15) (3, 7)
        8'b10101010, // Color (7, 15, 15) (4, 7)
        8'b10101010, // Color (7, 15, 15) (5, 7)
        8'b10101000, // Color (6, 15, 14) (6, 7)
        8'b10101000, // Color (6, 15, 14) (7, 7)
        8'b10101010, // Color (7, 15, 15) (8, 7)
        8'b10101010, // Color (7, 15, 15) (9, 7)
        8'b10101000, // Color (6, 15, 14) (10, 7)
        8'b10011110, // Color (4, 14, 14) (11, 7)
        8'b10011110, // Color (4, 14, 14) (12, 7)
        8'b10100000, // Color (3, 14, 14) (13, 7)
        8'b10011110, // Color (4, 14, 14) (14, 7)
        8'b10101100, // Color (0, 11, 11) (15, 7)
        8'b10100000, // Color (3, 14, 14) (0, 8)
        8'b10100110, // Color (9, 15, 14) (1, 8)
        8'b10101010, // Color (7, 15, 15) (2, 8)
        8'b10101010, // Color (7, 15, 15) (3, 8)
        8'b10101010, // Color (7, 15, 15) (4, 8)
        8'b10101000, // Color (6, 15, 14) (5, 8)
        8'b10101000, // Color (6, 15, 14) (6, 8)
        8'b10101010, // Color (7, 15, 15) (7, 8)
        8'b10101010, // Color (7, 15, 15) (8, 8)
        8'b10101000, // Color (6, 15, 14) (9, 8)
        8'b10101000, // Color (6, 15, 14) (10, 8)
        8'b10011110, // Color (4, 14, 14) (11, 8)
        8'b10011110, // Color (4, 14, 14) (12, 8)
        8'b10011110, // Color (4, 14, 14) (13, 8)
        8'b10101000, // Color (6, 15, 14) (14, 8)
        8'b10100010, // Color (1, 12, 12) (15, 8)
        8'b10100000, // Color (3, 14, 14) (0, 9)
        8'b10100110, // Color (9, 15, 14) (1, 9)
        8'b10101010, // Color (7, 15, 15) (2, 9)
        8'b10101010, // Color (7, 15, 15) (3, 9)
        8'b10101000, // Color (6, 15, 14) (4, 9)
        8'b10101000, // Color (6, 15, 14) (5, 9)
        8'b10101010, // Color (7, 15, 15) (6, 9)
        8'b10101010, // Color (7, 15, 15) (7, 9)
        8'b10101000, // Color (6, 15, 14) (8, 9)
        8'b10101000, // Color (6, 15, 14) (9, 9)
        8'b10101000, // Color (6, 15, 14) (10, 9)
        8'b10101000, // Color (6, 15, 14) (11, 9)
        8'b10011110, // Color (4, 14, 14) (12, 9)
        8'b10101010, // Color (7, 15, 15) (13, 9)
        8'b10101000, // Color (6, 15, 14) (14, 9)
        8'b10100010, // Color (1, 12, 12) (15, 9)
        8'b10100000, // Color (3, 14, 14) (0, 10)
        8'b10101000, // Color (6, 15, 14) (1, 10)
        8'b10101010, // Color (7, 15, 15) (2, 10)
        8'b10101000, // Color (6, 15, 14) (3, 10)
        8'b10101000, // Color (6, 15, 14) (4, 10)
        8'b10100110, // Color (9, 15, 14) (5, 10)
        8'b10100110, // Color (9, 15, 14) (6, 10)
        8'b10101000, // Color (6, 15, 14) (7, 10)
        8'b10101000, // Color (6, 15, 14) (8, 10)
        8'b10101000, // Color (6, 15, 14) (9, 10)
        8'b10101000, // Color (6, 15, 14) (10, 10)
        8'b10101000, // Color (6, 15, 14) (11, 10)
        8'b10100110, // Color (9, 15, 14) (12, 10)
        8'b10101010, // Color (7, 15, 15) (13, 10)
        8'b10011110, // Color (4, 14, 14) (14, 10)
        8'b10101100, // Color (0, 11, 11) (15, 10)
        8'b10100000, // Color (3, 14, 14) (0, 11)
        8'b10011110, // Color (4, 14, 14) (1, 11)
        8'b10101000, // Color (6, 15, 14) (2, 11)
        8'b10101000, // Color (6, 15, 14) (3, 11)
        8'b10100110, // Color (9, 15, 14) (4, 11)
        8'b10100110, // Color (9, 15, 14) (5, 11)
        8'b10101000, // Color (6, 15, 14) (6, 11)
        8'b10011110, // Color (4, 14, 14) (7, 11)
        8'b10011110, // Color (4, 14, 14) (8, 11)
        8'b10101000, // Color (6, 15, 14) (9, 11)
        8'b10011110, // Color (4, 14, 14) (10, 11)
        8'b10100110, // Color (9, 15, 14) (11, 11)
        8'b10100110, // Color (9, 15, 14) (12, 11)
        8'b10101000, // Color (6, 15, 14) (13, 11)
        8'b10011110, // Color (4, 14, 14) (14, 11)
        8'b10101100, // Color (0, 11, 11) (15, 11)
        8'b10100000, // Color (3, 14, 14) (0, 12)
        8'b10011110, // Color (4, 14, 14) (1, 12)
        8'b10101000, // Color (6, 15, 14) (2, 12)
        8'b10100110, // Color (9, 15, 14) (3, 12)
        8'b10100110, // Color (9, 15, 14) (4, 12)
        8'b10101000, // Color (6, 15, 14) (5, 12)
        8'b10011110, // Color (4, 14, 14) (6, 12)
        8'b10100000, // Color (3, 14, 14) (7, 12)
        8'b10100000, // Color (3, 14, 14) (8, 12)
        8'b10011110, // Color (4, 14, 14) (9, 12)
        8'b10101010, // Color (7, 15, 15) (10, 12)
        8'b10101010, // Color (7, 15, 15) (11, 12)
        8'b10101000, // Color (6, 15, 14) (12, 12)
        8'b10011110, // Color (4, 14, 14) (13, 12)
        8'b10101000, // Color (6, 15, 14) (14, 12)
        8'b10100010, // Color (1, 12, 12) (15, 12)
        8'b10100000, // Color (3, 14, 14) (0, 13)
        8'b10100000, // Color (3, 14, 14) (1, 13)
        8'b10101010, // Color (7, 15, 15) (2, 13)
        8'b10101010, // Color (7, 15, 15) (3, 13)
        8'b10101000, // Color (6, 15, 14) (4, 13)
        8'b10011110, // Color (4, 14, 14) (5, 13)
        8'b10100000, // Color (3, 14, 14) (6, 13)
        8'b10100000, // Color (3, 14, 14) (7, 13)
        8'b10011110, // Color (4, 14, 14) (8, 13)
        8'b10101000, // Color (6, 15, 14) (9, 13)
        8'b10101000, // Color (6, 15, 14) (10, 13)
        8'b10101000, // Color (6, 15, 14) (11, 13)
        8'b10011110, // Color (4, 14, 14) (12, 13)
        8'b10011110, // Color (4, 14, 14) (13, 13)
        8'b10101010, // Color (7, 15, 15) (14, 13)
        8'b10100010, // Color (1, 12, 12) (15, 13)
        8'b10100000, // Color (3, 14, 14) (0, 14)
        8'b10011110, // Color (4, 14, 14) (1, 14)
        8'b10100000, // Color (3, 14, 14) (2, 14)
        8'b10011110, // Color (4, 14, 14) (3, 14)
        8'b10011110, // Color (4, 14, 14) (4, 14)
        8'b10100000, // Color (3, 14, 14) (5, 14)
        8'b10100000, // Color (3, 14, 14) (6, 14)
        8'b10011110, // Color (4, 14, 14) (7, 14)
        8'b10101000, // Color (6, 15, 14) (8, 14)
        8'b10101000, // Color (6, 15, 14) (9, 14)
        8'b10011110, // Color (4, 14, 14) (10, 14)
        8'b10011110, // Color (4, 14, 14) (11, 14)
        8'b10101000, // Color (6, 15, 14) (12, 14)
        8'b10101010, // Color (7, 15, 15) (13, 14)
        8'b10100110, // Color (9, 15, 14) (14, 14)
        8'b10101100, // Color (0, 11, 11) (15, 14)
        8'b10100010, // Color (1, 12, 12) (0, 15)
        8'b10100010, // Color (1, 12, 12) (1, 15)
        8'b10101100, // Color (0, 11, 11) (2, 15)
        8'b10100010, // Color (1, 12, 12) (3, 15)
        8'b10100010, // Color (1, 12, 12) (4, 15)
        8'b10101100, // Color (0, 11, 11) (5, 15)
        8'b10101100, // Color (0, 11, 11) (6, 15)
        8'b10101100, // Color (0, 11, 11) (7, 15)
        8'b10100010, // Color (1, 12, 12) (8, 15)
        8'b10100010, // Color (1, 12, 12) (9, 15)
        8'b10101100, // Color (0, 11, 11) (10, 15)
        8'b10101100, // Color (0, 11, 11) (11, 15)
        8'b10100010, // Color (1, 12, 12) (12, 15)
        8'b10100010, // Color (1, 12, 12) (13, 15)
        8'b10101100, // Color (0, 11, 11) (14, 15)
        8'b10101100, // Color (0, 11, 11) (15, 15)
        // 18_furnace_front
        8'b10101110, // Color (5, 4, 4) (0, 0)
        8'b10101110, // Color (5, 4, 4) (1, 0)
        8'b10101110, // Color (5, 4, 4) (2, 0)
        8'b10101110, // Color (5, 4, 4) (3, 0)
        8'b10110000, // Color (3, 3, 3) (4, 0)
        8'b10101110, // Color (5, 4, 4) (5, 0)
        8'b10101110, // Color (5, 4, 4) (6, 0)
        8'b10101110, // Color (5, 4, 4) (7, 0)
        8'b10110000, // Color (3, 3, 3) (8, 0)
        8'b10110000, // Color (3, 3, 3) (9, 0)
        8'b10110000, // Color (3, 3, 3) (10, 0)
        8'b10101110, // Color (5, 4, 4) (11, 0)
        8'b10110000, // Color (3, 3, 3) (12, 0)
        8'b10110000, // Color (3, 3, 3) (13, 0)
        8'b10101110, // Color (5, 4, 4) (14, 0)
        8'b10101110, // Color (5, 4, 4) (15, 0)
        8'b10101110, // Color (5, 4, 4) (0, 1)
        8'b00001100, // Color (6, 6, 6) (1, 1)
        8'b00001100, // Color (6, 6, 6) (2, 1)
        8'b01011100, // Color (7, 7, 7) (3, 1)
        8'b01011100, // Color (7, 7, 7) (4, 1)
        8'b00001100, // Color (6, 6, 6) (5, 1)
        8'b01011100, // Color (7, 7, 7) (6, 1)
        8'b00001100, // Color (6, 6, 6) (7, 1)
        8'b01011100, // Color (7, 7, 7) (8, 1)
        8'b01011100, // Color (7, 7, 7) (9, 1)
        8'b00001100, // Color (6, 6, 6) (10, 1)
        8'b01011100, // Color (7, 7, 7) (11, 1)
        8'b00001100, // Color (6, 6, 6) (12, 1)
        8'b01011100, // Color (7, 7, 7) (13, 1)
        8'b01100100, // Color (5, 5, 5) (14, 1)
        8'b10101110, // Color (5, 4, 4) (15, 1)
        8'b10110000, // Color (3, 3, 3) (0, 2)
        8'b01100100, // Color (5, 5, 5) (1, 2)
        8'b01011100, // Color (7, 7, 7) (2, 2)
        8'b10110010, // Color (9, 9, 9) (3, 2)
        8'b01011100, // Color (7, 7, 7) (4, 2)
        8'b00001010, // Color (8, 8, 8) (5, 2)
        8'b00001100, // Color (6, 6, 6) (6, 2)
        8'b01011100, // Color (7, 7, 7) (7, 2)
        8'b00001010, // Color (8, 8, 8) (8, 2)
        8'b10110010, // Color (9, 9, 9) (9, 2)
        8'b00001010, // Color (8, 8, 8) (10, 2)
        8'b10110010, // Color (9, 9, 9) (11, 2)
        8'b01011100, // Color (7, 7, 7) (12, 2)
        8'b00001100, // Color (6, 6, 6) (13, 2)
        8'b01011100, // Color (7, 7, 7) (14, 2)
        8'b10101110, // Color (5, 4, 4) (15, 2)
        8'b10101110, // Color (5, 4, 4) (0, 3)
        8'b00001100, // Color (6, 6, 6) (1, 3)
        8'b00001010, // Color (8, 8, 8) (2, 3)
        8'b00001010, // Color (8, 8, 8) (3, 3)
        8'b10110000, // Color (3, 3, 3) (4, 3)
        8'b01010110, // Color (2, 2, 2) (5, 3)
        8'b01010110, // Color (2, 2, 2) (6, 3)
        8'b01010110, // Color (2, 2, 2) (7, 3)
        8'b01010110, // Color (2, 2, 2) (8, 3)
        8'b01010110, // Color (2, 2, 2) (9, 3)
        8'b01010110, // Color (2, 2, 2) (10, 3)
        8'b10110000, // Color (3, 3, 3) (11, 3)
        8'b00001010, // Color (8, 8, 8) (12, 3)
        8'b01011100, // Color (7, 7, 7) (13, 3)
        8'b00001100, // Color (6, 6, 6) (14, 3)
        8'b10101110, // Color (5, 4, 4) (15, 3)
        8'b10101110, // Color (5, 4, 4) (0, 4)
        8'b01011100, // Color (7, 7, 7) (1, 4)
        8'b00001010, // Color (8, 8, 8) (2, 4)
        8'b10110000, // Color (3, 3, 3) (3, 4)
        8'b01100000, // Color (1, 1, 1) (4, 4)
        8'b01100000, // Color (1, 1, 1) (5, 4)
        8'b01100000, // Color (1, 1, 1) (6, 4)
        8'b01100000, // Color (1, 1, 1) (7, 4)
        8'b01100000, // Color (1, 1, 1) (8, 4)
        8'b01100000, // Color (1, 1, 1) (9, 4)
        8'b01100000, // Color (1, 1, 1) (10, 4)
        8'b01100000, // Color (1, 1, 1) (11, 4)
        8'b10110000, // Color (3, 3, 3) (12, 4)
        8'b01011100, // Color (7, 7, 7) (13, 4)
        8'b01100100, // Color (5, 5, 5) (14, 4)
        8'b10110000, // Color (3, 3, 3) (15, 4)
        8'b10110000, // Color (3, 3, 3) (0, 5)
        8'b01011100, // Color (7, 7, 7) (1, 5)
        8'b00001100, // Color (6, 6, 6) (2, 5)
        8'b01100000, // Color (1, 1, 1) (3, 5)
        8'b01100000, // Color (1, 1, 1) (4, 5)
        8'b01100000, // Color (1, 1, 1) (5, 5)
        8'b01010110, // Color (2, 2, 2) (6, 5)
        8'b01010110, // Color (2, 2, 2) (7, 5)
        8'b01010110, // Color (2, 2, 2) (8, 5)
        8'b01010110, // Color (2, 2, 2) (9, 5)
        8'b01100000, // Color (1, 1, 1) (10, 5)
        8'b01100000, // Color (1, 1, 1) (11, 5)
        8'b01100000, // Color (1, 1, 1) (12, 5)
        8'b10110010, // Color (9, 9, 9) (13, 5)
        8'b01100100, // Color (5, 5, 5) (14, 5)
        8'b10110000, // Color (3, 3, 3) (15, 5)
        8'b10101110, // Color (5, 4, 4) (0, 6)
        8'b01011100, // Color (7, 7, 7) (1, 6)
        8'b00001100, // Color (6, 6, 6) (2, 6)
        8'b01100000, // Color (1, 1, 1) (3, 6)
        8'b01100000, // Color (1, 1, 1) (4, 6)
        8'b10110000, // Color (3, 3, 3) (5, 6)
        8'b10110000, // Color (3, 3, 3) (6, 6)
        8'b10110000, // Color (3, 3, 3) (7, 6)
        8'b10110000, // Color (3, 3, 3) (8, 6)
        8'b10110000, // Color (3, 3, 3) (9, 6)
        8'b10110000, // Color (3, 3, 3) (10, 6)
        8'b01100000, // Color (1, 1, 1) (11, 6)
        8'b01100000, // Color (1, 1, 1) (12, 6)
        8'b10110010, // Color (9, 9, 9) (13, 6)
        8'b01100100, // Color (5, 5, 5) (14, 6)
        8'b10101110, // Color (5, 4, 4) (15, 6)
        8'b10110000, // Color (3, 3, 3) (0, 7)
        8'b01011100, // Color (7, 7, 7) (1, 7)
        8'b10110010, // Color (9, 9, 9) (2, 7)
        8'b01100010, // Color (10, 10, 10) (3, 7)
        8'b01100010, // Color (10, 10, 10) (4, 7)
        8'b01100110, // Color (11, 11, 11) (5, 7)
        8'b01100110, // Color (11, 11, 11) (6, 7)
        8'b01100110, // Color (11, 11, 11) (7, 7)
        8'b01100110, // Color (11, 11, 11) (8, 7)
        8'b01100110, // Color (11, 11, 11) (9, 7)
        8'b01100110, // Color (11, 11, 11) (10, 7)
        8'b01100010, // Color (10, 10, 10) (11, 7)
        8'b01100010, // Color (10, 10, 10) (12, 7)
        8'b10110010, // Color (9, 9, 9) (13, 7)
        8'b01011100, // Color (7, 7, 7) (14, 7)
        8'b10110000, // Color (3, 3, 3) (15, 7)
        8'b10110000, // Color (3, 3, 3) (0, 8)
        8'b01011100, // Color (7, 7, 7) (1, 8)
        8'b00001010, // Color (8, 8, 8) (2, 8)
        8'b01011100, // Color (7, 7, 7) (3, 8)
        8'b00001100, // Color (6, 6, 6) (4, 8)
        8'b01100100, // Color (5, 5, 5) (5, 8)
        8'b01011100, // Color (7, 7, 7) (6, 8)
        8'b00001100, // Color (6, 6, 6) (7, 8)
        8'b01100100, // Color (5, 5, 5) (8, 8)
        8'b00001100, // Color (6, 6, 6) (9, 8)
        8'b01011100, // Color (7, 7, 7) (10, 8)
        8'b00001100, // Color (6, 6, 6) (11, 8)
        8'b01011100, // Color (7, 7, 7) (12, 8)
        8'b00001100, // Color (6, 6, 6) (13, 8)
        8'b00001100, // Color (6, 6, 6) (14, 8)
        8'b10101110, // Color (5, 4, 4) (15, 8)
        8'b10101110, // Color (5, 4, 4) (0, 9)
        8'b10000000, // Color (12, 12, 12) (1, 9)
        8'b01100110, // Color (11, 11, 11) (2, 9)
        8'b10000000, // Color (12, 12, 12) (3, 9)
        8'b10000000, // Color (12, 12, 12) (4, 9)
        8'b10000000, // Color (12, 12, 12) (5, 9)
        8'b10000000, // Color (12, 12, 12) (6, 9)
        8'b10000000, // Color (12, 12, 12) (7, 9)
        8'b10000000, // Color (12, 12, 12) (8, 9)
        8'b10000000, // Color (12, 12, 12) (9, 9)
        8'b10000000, // Color (12, 12, 12) (10, 9)
        8'b10000000, // Color (12, 12, 12) (11, 9)
        8'b10000000, // Color (12, 12, 12) (12, 9)
        8'b10000000, // Color (12, 12, 12) (13, 9)
        8'b01100010, // Color (10, 10, 10) (14, 9)
        8'b10101110, // Color (5, 4, 4) (15, 9)
        8'b10101110, // Color (5, 4, 4) (0, 10)
        8'b01100010, // Color (10, 10, 10) (1, 10)
        8'b01100010, // Color (10, 10, 10) (2, 10)
        8'b01100010, // Color (10, 10, 10) (3, 10)
        8'b01100110, // Color (11, 11, 11) (4, 10)
        8'b01100010, // Color (10, 10, 10) (5, 10)
        8'b00001010, // Color (8, 8, 8) (6, 10)
        8'b00001010, // Color (8, 8, 8) (7, 10)
        8'b00001010, // Color (8, 8, 8) (8, 10)
        8'b00001010, // Color (8, 8, 8) (9, 10)
        8'b01100010, // Color (10, 10, 10) (10, 10)
        8'b01100110, // Color (11, 11, 11) (11, 10)
        8'b01100010, // Color (10, 10, 10) (12, 10)
        8'b01100110, // Color (11, 11, 11) (13, 10)
        8'b10110010, // Color (9, 9, 9) (14, 10)
        8'b10110000, // Color (3, 3, 3) (15, 10)
        8'b10101110, // Color (5, 4, 4) (0, 11)
        8'b10110010, // Color (9, 9, 9) (1, 11)
        8'b01100010, // Color (10, 10, 10) (2, 11)
        8'b10110010, // Color (9, 9, 9) (3, 11)
        8'b01100100, // Color (5, 5, 5) (4, 11)
        8'b01010110, // Color (2, 2, 2) (5, 11)
        8'b01100000, // Color (1, 1, 1) (6, 11)
        8'b01100000, // Color (1, 1, 1) (7, 11)
        8'b01100000, // Color (1, 1, 1) (8, 11)
        8'b01100000, // Color (1, 1, 1) (9, 11)
        8'b01010110, // Color (2, 2, 2) (10, 11)
        8'b01100100, // Color (5, 5, 5) (11, 11)
        8'b10110010, // Color (9, 9, 9) (12, 11)
        8'b01100010, // Color (10, 10, 10) (13, 11)
        8'b10110010, // Color (9, 9, 9) (14, 11)
        8'b10101110, // Color (5, 4, 4) (15, 11)
        8'b10101110, // Color (5, 4, 4) (0, 12)
        8'b10110010, // Color (9, 9, 9) (1, 12)
        8'b10110010, // Color (9, 9, 9) (2, 12)
        8'b10101110, // Color (5, 4, 4) (3, 12)
        8'b01100000, // Color (1, 1, 1) (4, 12)
        8'b01100000, // Color (1, 1, 1) (5, 12)
        8'b01100000, // Color (1, 1, 1) (6, 12)
        8'b01100000, // Color (1, 1, 1) (7, 12)
        8'b01100000, // Color (1, 1, 1) (8, 12)
        8'b01100000, // Color (1, 1, 1) (9, 12)
        8'b01100000, // Color (1, 1, 1) (10, 12)
        8'b01100000, // Color (1, 1, 1) (11, 12)
        8'b10101110, // Color (5, 4, 4) (12, 12)
        8'b01011100, // Color (7, 7, 7) (13, 12)
        8'b10110010, // Color (9, 9, 9) (14, 12)
        8'b10101110, // Color (5, 4, 4) (15, 12)
        8'b10101110, // Color (5, 4, 4) (0, 13)
        8'b01011100, // Color (7, 7, 7) (1, 13)
        8'b10110010, // Color (9, 9, 9) (2, 13)
        8'b01100000, // Color (1, 1, 1) (3, 13)
        8'b01100000, // Color (1, 1, 1) (4, 13)
        8'b01100000, // Color (1, 1, 1) (5, 13)
        8'b01010110, // Color (2, 2, 2) (6, 13)
        8'b01010110, // Color (2, 2, 2) (7, 13)
        8'b01010110, // Color (2, 2, 2) (8, 13)
        8'b01010110, // Color (2, 2, 2) (9, 13)
        8'b01100000, // Color (1, 1, 1) (10, 13)
        8'b01100000, // Color (1, 1, 1) (11, 13)
        8'b01100000, // Color (1, 1, 1) (12, 13)
        8'b10110010, // Color (9, 9, 9) (13, 13)
        8'b10110010, // Color (9, 9, 9) (14, 13)
        8'b10101110, // Color (5, 4, 4) (15, 13)
        8'b10110000, // Color (3, 3, 3) (0, 14)
        8'b10110010, // Color (9, 9, 9) (1, 14)
        8'b01011100, // Color (7, 7, 7) (2, 14)
        8'b01100000, // Color (1, 1, 1) (3, 14)
        8'b01010110, // Color (2, 2, 2) (4, 14)
        8'b01010110, // Color (2, 2, 2) (5, 14)
        8'b01010110, // Color (2, 2, 2) (6, 14)
        8'b01010110, // Color (2, 2, 2) (7, 14)
        8'b01010110, // Color (2, 2, 2) (8, 14)
        8'b01010110, // Color (2, 2, 2) (9, 14)
        8'b01010110, // Color (2, 2, 2) (10, 14)
        8'b01010110, // Color (2, 2, 2) (11, 14)
        8'b01100000, // Color (1, 1, 1) (12, 14)
        8'b01011100, // Color (7, 7, 7) (13, 14)
        8'b10110010, // Color (9, 9, 9) (14, 14)
        8'b10110000, // Color (3, 3, 3) (15, 14)
        8'b10110000, // Color (3, 3, 3) (0, 15)
        8'b00001100, // Color (6, 6, 6) (1, 15)
        8'b10110000, // Color (3, 3, 3) (2, 15)
        8'b10110000, // Color (3, 3, 3) (3, 15)
        8'b10110000, // Color (3, 3, 3) (4, 15)
        8'b10101110, // Color (5, 4, 4) (5, 15)
        8'b10101110, // Color (5, 4, 4) (6, 15)
        8'b10101110, // Color (5, 4, 4) (7, 15)
        8'b10101110, // Color (5, 4, 4) (8, 15)
        8'b10101110, // Color (5, 4, 4) (9, 15)
        8'b10101110, // Color (5, 4, 4) (10, 15)
        8'b10110000, // Color (3, 3, 3) (11, 15)
        8'b10110000, // Color (3, 3, 3) (12, 15)
        8'b10110000, // Color (3, 3, 3) (13, 15)
        8'b00001100, // Color (6, 6, 6) (14, 15)
        8'b10110000, // Color (3, 3, 3) (15, 15)
        // 19_furnace_side
        8'b10101110, // Color (5, 4, 4) (0, 0)
        8'b10101110, // Color (5, 4, 4) (1, 0)
        8'b10101110, // Color (5, 4, 4) (2, 0)
        8'b10101110, // Color (5, 4, 4) (3, 0)
        8'b10110000, // Color (3, 3, 3) (4, 0)
        8'b10101110, // Color (5, 4, 4) (5, 0)
        8'b10101110, // Color (5, 4, 4) (6, 0)
        8'b10101110, // Color (5, 4, 4) (7, 0)
        8'b10110000, // Color (3, 3, 3) (8, 0)
        8'b10110000, // Color (3, 3, 3) (9, 0)
        8'b10110000, // Color (3, 3, 3) (10, 0)
        8'b10101110, // Color (5, 4, 4) (11, 0)
        8'b10110000, // Color (3, 3, 3) (12, 0)
        8'b10110000, // Color (3, 3, 3) (13, 0)
        8'b10101110, // Color (5, 4, 4) (14, 0)
        8'b10101110, // Color (5, 4, 4) (15, 0)
        8'b10101110, // Color (5, 4, 4) (0, 1)
        8'b01100100, // Color (5, 5, 5) (1, 1)
        8'b00001100, // Color (6, 6, 6) (2, 1)
        8'b00001100, // Color (6, 6, 6) (3, 1)
        8'b01011100, // Color (7, 7, 7) (4, 1)
        8'b00001100, // Color (6, 6, 6) (5, 1)
        8'b00001010, // Color (8, 8, 8) (6, 1)
        8'b01011100, // Color (7, 7, 7) (7, 1)
        8'b00001100, // Color (6, 6, 6) (8, 1)
        8'b00001100, // Color (6, 6, 6) (9, 1)
        8'b00001100, // Color (6, 6, 6) (10, 1)
        8'b01011100, // Color (7, 7, 7) (11, 1)
        8'b00001100, // Color (6, 6, 6) (12, 1)
        8'b00001100, // Color (6, 6, 6) (13, 1)
        8'b01100100, // Color (5, 5, 5) (14, 1)
        8'b10101110, // Color (5, 4, 4) (15, 1)
        8'b10101110, // Color (5, 4, 4) (0, 2)
        8'b01100100, // Color (5, 5, 5) (1, 2)
        8'b01011100, // Color (7, 7, 7) (2, 2)
        8'b10110010, // Color (9, 9, 9) (3, 2)
        8'b10110010, // Color (9, 9, 9) (4, 2)
        8'b01100100, // Color (5, 5, 5) (5, 2)
        8'b00001100, // Color (6, 6, 6) (6, 2)
        8'b01100100, // Color (5, 5, 5) (7, 2)
        8'b00001010, // Color (8, 8, 8) (8, 2)
        8'b00001010, // Color (8, 8, 8) (9, 2)
        8'b01011100, // Color (7, 7, 7) (10, 2)
        8'b00001100, // Color (6, 6, 6) (11, 2)
        8'b00001010, // Color (8, 8, 8) (12, 2)
        8'b00001010, // Color (8, 8, 8) (13, 2)
        8'b01011100, // Color (7, 7, 7) (14, 2)
        8'b10101110, // Color (5, 4, 4) (15, 2)
        8'b10101110, // Color (5, 4, 4) (0, 3)
        8'b00001100, // Color (6, 6, 6) (1, 3)
        8'b00001010, // Color (8, 8, 8) (2, 3)
        8'b00001010, // Color (8, 8, 8) (3, 3)
        8'b00001010, // Color (8, 8, 8) (4, 3)
        8'b10110010, // Color (9, 9, 9) (5, 3)
        8'b01100100, // Color (5, 5, 5) (6, 3)
        8'b00001100, // Color (6, 6, 6) (7, 3)
        8'b01011100, // Color (7, 7, 7) (8, 3)
        8'b10110010, // Color (9, 9, 9) (9, 3)
        8'b00001010, // Color (8, 8, 8) (10, 3)
        8'b00001010, // Color (8, 8, 8) (11, 3)
        8'b00001100, // Color (6, 6, 6) (12, 3)
        8'b00001010, // Color (8, 8, 8) (13, 3)
        8'b00001010, // Color (8, 8, 8) (14, 3)
        8'b10101110, // Color (5, 4, 4) (15, 3)
        8'b10101110, // Color (5, 4, 4) (0, 4)
        8'b01100100, // Color (5, 5, 5) (1, 4)
        8'b01011100, // Color (7, 7, 7) (2, 4)
        8'b00001010, // Color (8, 8, 8) (3, 4)
        8'b00001010, // Color (8, 8, 8) (4, 4)
        8'b01011100, // Color (7, 7, 7) (5, 4)
        8'b01100100, // Color (5, 5, 5) (6, 4)
        8'b01011100, // Color (7, 7, 7) (7, 4)
        8'b00001100, // Color (6, 6, 6) (8, 4)
        8'b00001010, // Color (8, 8, 8) (9, 4)
        8'b10110010, // Color (9, 9, 9) (10, 4)
        8'b00001010, // Color (8, 8, 8) (11, 4)
        8'b01100100, // Color (5, 5, 5) (12, 4)
        8'b01011100, // Color (7, 7, 7) (13, 4)
        8'b00001100, // Color (6, 6, 6) (14, 4)
        8'b10110000, // Color (3, 3, 3) (15, 4)
        8'b10110000, // Color (3, 3, 3) (0, 5)
        8'b01100100, // Color (5, 5, 5) (1, 5)
        8'b01100100, // Color (5, 5, 5) (2, 5)
        8'b00001100, // Color (6, 6, 6) (3, 5)
        8'b00001100, // Color (6, 6, 6) (4, 5)
        8'b01100100, // Color (5, 5, 5) (5, 5)
        8'b00001010, // Color (8, 8, 8) (6, 5)
        8'b10110010, // Color (9, 9, 9) (7, 5)
        8'b00001010, // Color (8, 8, 8) (8, 5)
        8'b00001100, // Color (6, 6, 6) (9, 5)
        8'b01011100, // Color (7, 7, 7) (10, 5)
        8'b00001010, // Color (8, 8, 8) (11, 5)
        8'b00001100, // Color (6, 6, 6) (12, 5)
        8'b10101110, // Color (5, 4, 4) (13, 5)
        8'b10101110, // Color (5, 4, 4) (14, 5)
        8'b10110000, // Color (3, 3, 3) (15, 5)
        8'b10101110, // Color (5, 4, 4) (0, 6)
        8'b00001100, // Color (6, 6, 6) (1, 6)
        8'b10110010, // Color (9, 9, 9) (2, 6)
        8'b10110010, // Color (9, 9, 9) (3, 6)
        8'b01011100, // Color (7, 7, 7) (4, 6)
        8'b00001100, // Color (6, 6, 6) (5, 6)
        8'b00001010, // Color (8, 8, 8) (6, 6)
        8'b00001010, // Color (8, 8, 8) (7, 6)
        8'b10110010, // Color (9, 9, 9) (8, 6)
        8'b00001010, // Color (8, 8, 8) (9, 6)
        8'b00001100, // Color (6, 6, 6) (10, 6)
        8'b00001100, // Color (6, 6, 6) (11, 6)
        8'b01011100, // Color (7, 7, 7) (12, 6)
        8'b01011100, // Color (7, 7, 7) (13, 6)
        8'b01100100, // Color (5, 5, 5) (14, 6)
        8'b10101110, // Color (5, 4, 4) (15, 6)
        8'b10110000, // Color (3, 3, 3) (0, 7)
        8'b01011100, // Color (7, 7, 7) (1, 7)
        8'b00001010, // Color (8, 8, 8) (2, 7)
        8'b00001010, // Color (8, 8, 8) (3, 7)
        8'b10110010, // Color (9, 9, 9) (4, 7)
        8'b00001100, // Color (6, 6, 6) (5, 7)
        8'b00001010, // Color (8, 8, 8) (6, 7)
        8'b00001010, // Color (8, 8, 8) (7, 7)
        8'b01011100, // Color (7, 7, 7) (8, 7)
        8'b01100100, // Color (5, 5, 5) (9, 7)
        8'b10110010, // Color (9, 9, 9) (10, 7)
        8'b00001010, // Color (8, 8, 8) (11, 7)
        8'b00001010, // Color (8, 8, 8) (12, 7)
        8'b00001010, // Color (8, 8, 8) (13, 7)
        8'b01011100, // Color (7, 7, 7) (14, 7)
        8'b10110000, // Color (3, 3, 3) (15, 7)
        8'b10110000, // Color (3, 3, 3) (0, 8)
        8'b00001100, // Color (6, 6, 6) (1, 8)
        8'b01011100, // Color (7, 7, 7) (2, 8)
        8'b01011100, // Color (7, 7, 7) (3, 8)
        8'b00001100, // Color (6, 6, 6) (4, 8)
        8'b01100100, // Color (5, 5, 5) (5, 8)
        8'b01100100, // Color (5, 5, 5) (6, 8)
        8'b01011100, // Color (7, 7, 7) (7, 8)
        8'b01100100, // Color (5, 5, 5) (8, 8)
        8'b10110010, // Color (9, 9, 9) (9, 8)
        8'b00001010, // Color (8, 8, 8) (10, 8)
        8'b00001010, // Color (8, 8, 8) (11, 8)
        8'b00001010, // Color (8, 8, 8) (12, 8)
        8'b01011100, // Color (7, 7, 7) (13, 8)
        8'b00001100, // Color (6, 6, 6) (14, 8)
        8'b10101110, // Color (5, 4, 4) (15, 8)
        8'b10101110, // Color (5, 4, 4) (0, 9)
        8'b10000000, // Color (12, 12, 12) (1, 9)
        8'b01100110, // Color (11, 11, 11) (2, 9)
        8'b10000000, // Color (12, 12, 12) (3, 9)
        8'b10000000, // Color (12, 12, 12) (4, 9)
        8'b10000000, // Color (12, 12, 12) (5, 9)
        8'b10000000, // Color (12, 12, 12) (6, 9)
        8'b10000000, // Color (12, 12, 12) (7, 9)
        8'b10000000, // Color (12, 12, 12) (8, 9)
        8'b10000000, // Color (12, 12, 12) (9, 9)
        8'b10000000, // Color (12, 12, 12) (10, 9)
        8'b10000000, // Color (12, 12, 12) (11, 9)
        8'b10000000, // Color (12, 12, 12) (12, 9)
        8'b10000000, // Color (12, 12, 12) (13, 9)
        8'b01100010, // Color (10, 10, 10) (14, 9)
        8'b10101110, // Color (5, 4, 4) (15, 9)
        8'b10101110, // Color (5, 4, 4) (0, 10)
        8'b10110010, // Color (9, 9, 9) (1, 10)
        8'b01100010, // Color (10, 10, 10) (2, 10)
        8'b01100010, // Color (10, 10, 10) (3, 10)
        8'b01100110, // Color (11, 11, 11) (4, 10)
        8'b01100010, // Color (10, 10, 10) (5, 10)
        8'b01100110, // Color (11, 11, 11) (6, 10)
        8'b01100110, // Color (11, 11, 11) (7, 10)
        8'b01100110, // Color (11, 11, 11) (8, 10)
        8'b01100110, // Color (11, 11, 11) (9, 10)
        8'b01100110, // Color (11, 11, 11) (10, 10)
        8'b01100110, // Color (11, 11, 11) (11, 10)
        8'b10110010, // Color (9, 9, 9) (12, 10)
        8'b01100110, // Color (11, 11, 11) (13, 10)
        8'b10110010, // Color (9, 9, 9) (14, 10)
        8'b10110000, // Color (3, 3, 3) (15, 10)
        8'b10110000, // Color (3, 3, 3) (0, 11)
        8'b10110010, // Color (9, 9, 9) (1, 11)
        8'b10110010, // Color (9, 9, 9) (2, 11)
        8'b01100010, // Color (10, 10, 10) (3, 11)
        8'b01100010, // Color (10, 10, 10) (4, 11)
        8'b01100010, // Color (10, 10, 10) (5, 11)
        8'b01100010, // Color (10, 10, 10) (6, 11)
        8'b01100010, // Color (10, 10, 10) (7, 11)
        8'b01100010, // Color (10, 10, 10) (8, 11)
        8'b01100010, // Color (10, 10, 10) (9, 11)
        8'b01100010, // Color (10, 10, 10) (10, 11)
        8'b01100010, // Color (10, 10, 10) (11, 11)
        8'b01100010, // Color (10, 10, 10) (12, 11)
        8'b01100010, // Color (10, 10, 10) (13, 11)
        8'b10110010, // Color (9, 9, 9) (14, 11)
        8'b10101110, // Color (5, 4, 4) (15, 11)
        8'b10110000, // Color (3, 3, 3) (0, 12)
        8'b10110010, // Color (9, 9, 9) (1, 12)
        8'b10110010, // Color (9, 9, 9) (2, 12)
        8'b10110010, // Color (9, 9, 9) (3, 12)
        8'b10110010, // Color (9, 9, 9) (4, 12)
        8'b10110010, // Color (9, 9, 9) (5, 12)
        8'b01100010, // Color (10, 10, 10) (6, 12)
        8'b10110010, // Color (9, 9, 9) (7, 12)
        8'b01100010, // Color (10, 10, 10) (8, 12)
        8'b01100010, // Color (10, 10, 10) (9, 12)
        8'b01100010, // Color (10, 10, 10) (10, 12)
        8'b01100010, // Color (10, 10, 10) (11, 12)
        8'b01100010, // Color (10, 10, 10) (12, 12)
        8'b10110010, // Color (9, 9, 9) (13, 12)
        8'b10110010, // Color (9, 9, 9) (14, 12)
        8'b10101110, // Color (5, 4, 4) (15, 12)
        8'b10101110, // Color (5, 4, 4) (0, 13)
        8'b01011100, // Color (7, 7, 7) (1, 13)
        8'b10110010, // Color (9, 9, 9) (2, 13)
        8'b10110010, // Color (9, 9, 9) (3, 13)
        8'b10110010, // Color (9, 9, 9) (4, 13)
        8'b10110010, // Color (9, 9, 9) (5, 13)
        8'b10110010, // Color (9, 9, 9) (6, 13)
        8'b10110010, // Color (9, 9, 9) (7, 13)
        8'b10110010, // Color (9, 9, 9) (8, 13)
        8'b01100010, // Color (10, 10, 10) (9, 13)
        8'b10110010, // Color (9, 9, 9) (10, 13)
        8'b10110010, // Color (9, 9, 9) (11, 13)
        8'b10110010, // Color (9, 9, 9) (12, 13)
        8'b10110010, // Color (9, 9, 9) (13, 13)
        8'b01011100, // Color (7, 7, 7) (14, 13)
        8'b10101110, // Color (5, 4, 4) (15, 13)
        8'b10101110, // Color (5, 4, 4) (0, 14)
        8'b00001100, // Color (6, 6, 6) (1, 14)
        8'b00001100, // Color (6, 6, 6) (2, 14)
        8'b01011100, // Color (7, 7, 7) (3, 14)
        8'b01011100, // Color (7, 7, 7) (4, 14)
        8'b00001100, // Color (6, 6, 6) (5, 14)
        8'b01011100, // Color (7, 7, 7) (6, 14)
        8'b01011100, // Color (7, 7, 7) (7, 14)
        8'b01011100, // Color (7, 7, 7) (8, 14)
        8'b01011100, // Color (7, 7, 7) (9, 14)
        8'b01011100, // Color (7, 7, 7) (10, 14)
        8'b01011100, // Color (7, 7, 7) (11, 14)
        8'b00001100, // Color (6, 6, 6) (12, 14)
        8'b00001100, // Color (6, 6, 6) (13, 14)
        8'b00001100, // Color (6, 6, 6) (14, 14)
        8'b10101110, // Color (5, 4, 4) (15, 14)
        8'b10101110, // Color (5, 4, 4) (0, 15)
        8'b10101110, // Color (5, 4, 4) (1, 15)
        8'b10101110, // Color (5, 4, 4) (2, 15)
        8'b10101110, // Color (5, 4, 4) (3, 15)
        8'b10110000, // Color (3, 3, 3) (4, 15)
        8'b10101110, // Color (5, 4, 4) (5, 15)
        8'b10101110, // Color (5, 4, 4) (6, 15)
        8'b10101110, // Color (5, 4, 4) (7, 15)
        8'b10110000, // Color (3, 3, 3) (8, 15)
        8'b10110000, // Color (3, 3, 3) (9, 15)
        8'b10110000, // Color (3, 3, 3) (10, 15)
        8'b10110000, // Color (3, 3, 3) (11, 15)
        8'b10101110, // Color (5, 4, 4) (12, 15)
        8'b10101110, // Color (5, 4, 4) (13, 15)
        8'b10101110, // Color (5, 4, 4) (14, 15)
        8'b10101110, // Color (5, 4, 4) (15, 15)
        // 20_furnace_top
        8'b10101110, // Color (5, 4, 4) (0, 0)
        8'b10101110, // Color (5, 4, 4) (1, 0)
        8'b10101110, // Color (5, 4, 4) (2, 0)
        8'b10101110, // Color (5, 4, 4) (3, 0)
        8'b10110000, // Color (3, 3, 3) (4, 0)
        8'b10101110, // Color (5, 4, 4) (5, 0)
        8'b10101110, // Color (5, 4, 4) (6, 0)
        8'b10101110, // Color (5, 4, 4) (7, 0)
        8'b10110000, // Color (3, 3, 3) (8, 0)
        8'b10110000, // Color (3, 3, 3) (9, 0)
        8'b10110000, // Color (3, 3, 3) (10, 0)
        8'b10101110, // Color (5, 4, 4) (11, 0)
        8'b10110000, // Color (3, 3, 3) (12, 0)
        8'b10110000, // Color (3, 3, 3) (13, 0)
        8'b10101110, // Color (5, 4, 4) (14, 0)
        8'b10101110, // Color (5, 4, 4) (15, 0)
        8'b10101110, // Color (5, 4, 4) (0, 1)
        8'b01100100, // Color (5, 5, 5) (1, 1)
        8'b01100100, // Color (5, 5, 5) (2, 1)
        8'b01100100, // Color (5, 5, 5) (3, 1)
        8'b00001100, // Color (6, 6, 6) (4, 1)
        8'b00001010, // Color (8, 8, 8) (5, 1)
        8'b00001010, // Color (8, 8, 8) (6, 1)
        8'b01011100, // Color (7, 7, 7) (7, 1)
        8'b01100100, // Color (5, 5, 5) (8, 1)
        8'b00001100, // Color (6, 6, 6) (9, 1)
        8'b00001100, // Color (6, 6, 6) (10, 1)
        8'b01011100, // Color (7, 7, 7) (11, 1)
        8'b00001010, // Color (8, 8, 8) (12, 1)
        8'b00001100, // Color (6, 6, 6) (13, 1)
        8'b01100100, // Color (5, 5, 5) (14, 1)
        8'b10101110, // Color (5, 4, 4) (15, 1)
        8'b10101110, // Color (5, 4, 4) (0, 2)
        8'b01100100, // Color (5, 5, 5) (1, 2)
        8'b01011100, // Color (7, 7, 7) (2, 2)
        8'b10110010, // Color (9, 9, 9) (3, 2)
        8'b10110010, // Color (9, 9, 9) (4, 2)
        8'b01011100, // Color (7, 7, 7) (5, 2)
        8'b01011100, // Color (7, 7, 7) (6, 2)
        8'b01100100, // Color (5, 5, 5) (7, 2)
        8'b00001010, // Color (8, 8, 8) (8, 2)
        8'b10110010, // Color (9, 9, 9) (9, 2)
        8'b00001010, // Color (8, 8, 8) (10, 2)
        8'b00001100, // Color (6, 6, 6) (11, 2)
        8'b00001010, // Color (8, 8, 8) (12, 2)
        8'b00001010, // Color (8, 8, 8) (13, 2)
        8'b01011100, // Color (7, 7, 7) (14, 2)
        8'b10101110, // Color (5, 4, 4) (15, 2)
        8'b10101110, // Color (5, 4, 4) (0, 3)
        8'b00001100, // Color (6, 6, 6) (1, 3)
        8'b10110010, // Color (9, 9, 9) (2, 3)
        8'b00001010, // Color (8, 8, 8) (3, 3)
        8'b10110010, // Color (9, 9, 9) (4, 3)
        8'b10110010, // Color (9, 9, 9) (5, 3)
        8'b01100100, // Color (5, 5, 5) (6, 3)
        8'b01011100, // Color (7, 7, 7) (7, 3)
        8'b10110010, // Color (9, 9, 9) (8, 3)
        8'b10110010, // Color (9, 9, 9) (9, 3)
        8'b10110010, // Color (9, 9, 9) (10, 3)
        8'b00001010, // Color (8, 8, 8) (11, 3)
        8'b00001100, // Color (6, 6, 6) (12, 3)
        8'b01011100, // Color (7, 7, 7) (13, 3)
        8'b01011100, // Color (7, 7, 7) (14, 3)
        8'b10101110, // Color (5, 4, 4) (15, 3)
        8'b10101110, // Color (5, 4, 4) (0, 4)
        8'b01011100, // Color (7, 7, 7) (1, 4)
        8'b00001010, // Color (8, 8, 8) (2, 4)
        8'b10110010, // Color (9, 9, 9) (3, 4)
        8'b00001010, // Color (8, 8, 8) (4, 4)
        8'b01011100, // Color (7, 7, 7) (5, 4)
        8'b01100100, // Color (5, 5, 5) (6, 4)
        8'b00001100, // Color (6, 6, 6) (7, 4)
        8'b01011100, // Color (7, 7, 7) (8, 4)
        8'b10110010, // Color (9, 9, 9) (9, 4)
        8'b10110010, // Color (9, 9, 9) (10, 4)
        8'b10110010, // Color (9, 9, 9) (11, 4)
        8'b01100100, // Color (5, 5, 5) (12, 4)
        8'b01011100, // Color (7, 7, 7) (13, 4)
        8'b00001100, // Color (6, 6, 6) (14, 4)
        8'b10110000, // Color (3, 3, 3) (15, 4)
        8'b10110000, // Color (3, 3, 3) (0, 5)
        8'b00001100, // Color (6, 6, 6) (1, 5)
        8'b01100100, // Color (5, 5, 5) (2, 5)
        8'b00001100, // Color (6, 6, 6) (3, 5)
        8'b00001100, // Color (6, 6, 6) (4, 5)
        8'b01100100, // Color (5, 5, 5) (5, 5)
        8'b00001010, // Color (8, 8, 8) (6, 5)
        8'b01011100, // Color (7, 7, 7) (7, 5)
        8'b00001100, // Color (6, 6, 6) (8, 5)
        8'b00001100, // Color (6, 6, 6) (9, 5)
        8'b01011100, // Color (7, 7, 7) (10, 5)
        8'b00001010, // Color (8, 8, 8) (11, 5)
        8'b01100100, // Color (5, 5, 5) (12, 5)
        8'b01100100, // Color (5, 5, 5) (13, 5)
        8'b10101110, // Color (5, 4, 4) (14, 5)
        8'b10110000, // Color (3, 3, 3) (15, 5)
        8'b10101110, // Color (5, 4, 4) (0, 6)
        8'b01100100, // Color (5, 5, 5) (1, 6)
        8'b00001010, // Color (8, 8, 8) (2, 6)
        8'b10110010, // Color (9, 9, 9) (3, 6)
        8'b00001100, // Color (6, 6, 6) (4, 6)
        8'b00001010, // Color (8, 8, 8) (5, 6)
        8'b10110010, // Color (9, 9, 9) (6, 6)
        8'b10110010, // Color (9, 9, 9) (7, 6)
        8'b10110010, // Color (9, 9, 9) (8, 6)
        8'b00001010, // Color (8, 8, 8) (9, 6)
        8'b01100100, // Color (5, 5, 5) (10, 6)
        8'b01100100, // Color (5, 5, 5) (11, 6)
        8'b00001010, // Color (8, 8, 8) (12, 6)
        8'b00001010, // Color (8, 8, 8) (13, 6)
        8'b00001100, // Color (6, 6, 6) (14, 6)
        8'b10101110, // Color (5, 4, 4) (15, 6)
        8'b10110000, // Color (3, 3, 3) (0, 7)
        8'b01011100, // Color (7, 7, 7) (1, 7)
        8'b10110010, // Color (9, 9, 9) (2, 7)
        8'b10110010, // Color (9, 9, 9) (3, 7)
        8'b00001010, // Color (8, 8, 8) (4, 7)
        8'b00001100, // Color (6, 6, 6) (5, 7)
        8'b10110010, // Color (9, 9, 9) (6, 7)
        8'b10110010, // Color (9, 9, 9) (7, 7)
        8'b10110010, // Color (9, 9, 9) (8, 7)
        8'b00001100, // Color (6, 6, 6) (9, 7)
        8'b00001010, // Color (8, 8, 8) (10, 7)
        8'b10110010, // Color (9, 9, 9) (11, 7)
        8'b10110010, // Color (9, 9, 9) (12, 7)
        8'b10110010, // Color (9, 9, 9) (13, 7)
        8'b01011100, // Color (7, 7, 7) (14, 7)
        8'b10110000, // Color (3, 3, 3) (15, 7)
        8'b10110000, // Color (3, 3, 3) (0, 8)
        8'b10110010, // Color (9, 9, 9) (1, 8)
        8'b10110010, // Color (9, 9, 9) (2, 8)
        8'b10110010, // Color (9, 9, 9) (3, 8)
        8'b10110010, // Color (9, 9, 9) (4, 8)
        8'b01011100, // Color (7, 7, 7) (5, 8)
        8'b01011100, // Color (7, 7, 7) (6, 8)
        8'b00001010, // Color (8, 8, 8) (7, 8)
        8'b00001100, // Color (6, 6, 6) (8, 8)
        8'b00001010, // Color (8, 8, 8) (9, 8)
        8'b10110010, // Color (9, 9, 9) (10, 8)
        8'b10110010, // Color (9, 9, 9) (11, 8)
        8'b10110010, // Color (9, 9, 9) (12, 8)
        8'b01011100, // Color (7, 7, 7) (13, 8)
        8'b00001010, // Color (8, 8, 8) (14, 8)
        8'b10101110, // Color (5, 4, 4) (15, 8)
        8'b10101110, // Color (5, 4, 4) (0, 9)
        8'b10110010, // Color (9, 9, 9) (1, 9)
        8'b10110010, // Color (9, 9, 9) (2, 9)
        8'b10110010, // Color (9, 9, 9) (3, 9)
        8'b10110010, // Color (9, 9, 9) (4, 9)
        8'b00001010, // Color (8, 8, 8) (5, 9)
        8'b00001100, // Color (6, 6, 6) (6, 9)
        8'b00001100, // Color (6, 6, 6) (7, 9)
        8'b00001010, // Color (8, 8, 8) (8, 9)
        8'b00001100, // Color (6, 6, 6) (9, 9)
        8'b01011100, // Color (7, 7, 7) (10, 9)
        8'b00001010, // Color (8, 8, 8) (11, 9)
        8'b00001010, // Color (8, 8, 8) (12, 9)
        8'b00001010, // Color (8, 8, 8) (13, 9)
        8'b10101110, // Color (5, 4, 4) (14, 9)
        8'b10101110, // Color (5, 4, 4) (15, 9)
        8'b10101110, // Color (5, 4, 4) (0, 10)
        8'b01011100, // Color (7, 7, 7) (1, 10)
        8'b10110010, // Color (9, 9, 9) (2, 10)
        8'b10110010, // Color (9, 9, 9) (3, 10)
        8'b10110010, // Color (9, 9, 9) (4, 10)
        8'b01011100, // Color (7, 7, 7) (5, 10)
        8'b00001010, // Color (8, 8, 8) (6, 10)
        8'b10110010, // Color (9, 9, 9) (7, 10)
        8'b10110010, // Color (9, 9, 9) (8, 10)
        8'b10110010, // Color (9, 9, 9) (9, 10)
        8'b00001010, // Color (8, 8, 8) (10, 10)
        8'b00001100, // Color (6, 6, 6) (11, 10)
        8'b01100100, // Color (5, 5, 5) (12, 10)
        8'b01100100, // Color (5, 5, 5) (13, 10)
        8'b00001100, // Color (6, 6, 6) (14, 10)
        8'b10110000, // Color (3, 3, 3) (15, 10)
        8'b10110000, // Color (3, 3, 3) (0, 11)
        8'b01100100, // Color (5, 5, 5) (1, 11)
        8'b01011100, // Color (7, 7, 7) (2, 11)
        8'b00001010, // Color (8, 8, 8) (3, 11)
        8'b01011100, // Color (7, 7, 7) (4, 11)
        8'b00001100, // Color (6, 6, 6) (5, 11)
        8'b10110010, // Color (9, 9, 9) (6, 11)
        8'b10110010, // Color (9, 9, 9) (7, 11)
        8'b10110010, // Color (9, 9, 9) (8, 11)
        8'b10110010, // Color (9, 9, 9) (9, 11)
        8'b10110010, // Color (9, 9, 9) (10, 11)
        8'b00001010, // Color (8, 8, 8) (11, 11)
        8'b00001100, // Color (6, 6, 6) (12, 11)
        8'b10110010, // Color (9, 9, 9) (13, 11)
        8'b01011100, // Color (7, 7, 7) (14, 11)
        8'b10101110, // Color (5, 4, 4) (15, 11)
        8'b10110000, // Color (3, 3, 3) (0, 12)
        8'b00001010, // Color (8, 8, 8) (1, 12)
        8'b01100100, // Color (5, 5, 5) (2, 12)
        8'b01100100, // Color (5, 5, 5) (3, 12)
        8'b00001100, // Color (6, 6, 6) (4, 12)
        8'b01100100, // Color (5, 5, 5) (5, 12)
        8'b01011100, // Color (7, 7, 7) (6, 12)
        8'b00001010, // Color (8, 8, 8) (7, 12)
        8'b10110010, // Color (9, 9, 9) (8, 12)
        8'b10110010, // Color (9, 9, 9) (9, 12)
        8'b10110010, // Color (9, 9, 9) (10, 12)
        8'b01011100, // Color (7, 7, 7) (11, 12)
        8'b00001010, // Color (8, 8, 8) (12, 12)
        8'b00001010, // Color (8, 8, 8) (13, 12)
        8'b00001010, // Color (8, 8, 8) (14, 12)
        8'b10101110, // Color (5, 4, 4) (15, 12)
        8'b10101110, // Color (5, 4, 4) (0, 13)
        8'b01011100, // Color (7, 7, 7) (1, 13)
        8'b10110010, // Color (9, 9, 9) (2, 13)
        8'b01100100, // Color (5, 5, 5) (3, 13)
        8'b01100100, // Color (5, 5, 5) (4, 13)
        8'b01011100, // Color (7, 7, 7) (5, 13)
        8'b01100100, // Color (5, 5, 5) (6, 13)
        8'b00001100, // Color (6, 6, 6) (7, 13)
        8'b01011100, // Color (7, 7, 7) (8, 13)
        8'b01011100, // Color (7, 7, 7) (9, 13)
        8'b01011100, // Color (7, 7, 7) (10, 13)
        8'b00001100, // Color (6, 6, 6) (11, 13)
        8'b00001010, // Color (8, 8, 8) (12, 13)
        8'b00001010, // Color (8, 8, 8) (13, 13)
        8'b01011100, // Color (7, 7, 7) (14, 13)
        8'b10101110, // Color (5, 4, 4) (15, 13)
        8'b10101110, // Color (5, 4, 4) (0, 14)
        8'b01100100, // Color (5, 5, 5) (1, 14)
        8'b01011100, // Color (7, 7, 7) (2, 14)
        8'b00001100, // Color (6, 6, 6) (3, 14)
        8'b01011100, // Color (7, 7, 7) (4, 14)
        8'b00001010, // Color (8, 8, 8) (5, 14)
        8'b01011100, // Color (7, 7, 7) (6, 14)
        8'b10101110, // Color (5, 4, 4) (7, 14)
        8'b01100100, // Color (5, 5, 5) (8, 14)
        8'b00001100, // Color (6, 6, 6) (9, 14)
        8'b00001100, // Color (6, 6, 6) (10, 14)
        8'b01100100, // Color (5, 5, 5) (11, 14)
        8'b00001100, // Color (6, 6, 6) (12, 14)
        8'b01011100, // Color (7, 7, 7) (13, 14)
        8'b00001100, // Color (6, 6, 6) (14, 14)
        8'b10101110, // Color (5, 4, 4) (15, 14)
        8'b10101110, // Color (5, 4, 4) (0, 15)
        8'b10101110, // Color (5, 4, 4) (1, 15)
        8'b10101110, // Color (5, 4, 4) (2, 15)
        8'b10101110, // Color (5, 4, 4) (3, 15)
        8'b10110000, // Color (3, 3, 3) (4, 15)
        8'b10101110, // Color (5, 4, 4) (5, 15)
        8'b10101110, // Color (5, 4, 4) (6, 15)
        8'b10101110, // Color (5, 4, 4) (7, 15)
        8'b10110000, // Color (3, 3, 3) (8, 15)
        8'b10110000, // Color (3, 3, 3) (9, 15)
        8'b10110000, // Color (3, 3, 3) (10, 15)
        8'b10110000, // Color (3, 3, 3) (11, 15)
        8'b10101110, // Color (5, 4, 4) (12, 15)
        8'b10101110, // Color (5, 4, 4) (13, 15)
        8'b10101110, // Color (5, 4, 4) (14, 15)
        8'b10101110, // Color (5, 4, 4) (15, 15)
        // 21_amethyst_block
        8'b10110100, // Color (6, 4, 9) (0, 0)
        8'b10110110, // Color (7, 5, 11) (1, 0)
        8'b10111000, // Color (8, 6, 12) (2, 0)
        8'b10110110, // Color (7, 5, 11) (3, 0)
        8'b10110110, // Color (7, 5, 11) (4, 0)
        8'b10110100, // Color (6, 4, 9) (5, 0)
        8'b10110110, // Color (7, 5, 11) (6, 0)
        8'b10111010, // Color (12, 9, 15) (7, 0)
        8'b10111100, // Color (15, 12, 14) (8, 0)
        8'b10111100, // Color (15, 12, 14) (9, 0)
        8'b10111110, // Color (10, 7, 15) (10, 0)
        8'b10111000, // Color (8, 6, 12) (11, 0)
        8'b10110100, // Color (6, 4, 9) (12, 0)
        8'b10110110, // Color (7, 5, 11) (13, 0)
        8'b10111000, // Color (8, 6, 12) (14, 0)
        8'b11000000, // Color (5, 3, 9) (15, 0)
        8'b10110110, // Color (7, 5, 11) (0, 1)
        8'b10111000, // Color (8, 6, 12) (1, 1)
        8'b10111110, // Color (10, 7, 15) (2, 1)
        8'b10111000, // Color (8, 6, 12) (3, 1)
        8'b10110100, // Color (6, 4, 9) (4, 1)
        8'b10110110, // Color (7, 5, 11) (5, 1)
        8'b10111000, // Color (8, 6, 12) (6, 1)
        8'b10110110, // Color (7, 5, 11) (7, 1)
        8'b10111000, // Color (8, 6, 12) (8, 1)
        8'b10111110, // Color (10, 7, 15) (9, 1)
        8'b11000000, // Color (5, 3, 9) (10, 1)
        8'b11000000, // Color (5, 3, 9) (11, 1)
        8'b10110110, // Color (7, 5, 11) (12, 1)
        8'b10111000, // Color (8, 6, 12) (13, 1)
        8'b10111000, // Color (8, 6, 12) (14, 1)
        8'b10110100, // Color (6, 4, 9) (15, 1)
        8'b10110100, // Color (6, 4, 9) (0, 2)
        8'b10111000, // Color (8, 6, 12) (1, 2)
        8'b10110110, // Color (7, 5, 11) (2, 2)
        8'b10110100, // Color (6, 4, 9) (3, 2)
        8'b10110100, // Color (6, 4, 9) (4, 2)
        8'b10111000, // Color (8, 6, 12) (5, 2)
        8'b10111110, // Color (10, 7, 15) (6, 2)
        8'b10110110, // Color (7, 5, 11) (7, 2)
        8'b10110100, // Color (6, 4, 9) (8, 2)
        8'b10111110, // Color (10, 7, 15) (9, 2)
        8'b11000000, // Color (5, 3, 9) (10, 2)
        8'b10110100, // Color (6, 4, 9) (11, 2)
        8'b10111110, // Color (10, 7, 15) (12, 2)
        8'b10110110, // Color (7, 5, 11) (13, 2)
        8'b10110110, // Color (7, 5, 11) (14, 2)
        8'b10110100, // Color (6, 4, 9) (15, 2)
        8'b10110100, // Color (6, 4, 9) (0, 3)
        8'b10110110, // Color (7, 5, 11) (1, 3)
        8'b10111000, // Color (8, 6, 12) (2, 3)
        8'b10110100, // Color (6, 4, 9) (3, 3)
        8'b11000000, // Color (5, 3, 9) (4, 3)
        8'b11000000, // Color (5, 3, 9) (5, 3)
        8'b10110110, // Color (7, 5, 11) (6, 3)
        8'b10110100, // Color (6, 4, 9) (7, 3)
        8'b10110100, // Color (6, 4, 9) (8, 3)
        8'b10110110, // Color (7, 5, 11) (9, 3)
        8'b10110100, // Color (6, 4, 9) (10, 3)
        8'b10111110, // Color (10, 7, 15) (11, 3)
        8'b10111010, // Color (12, 9, 15) (12, 3)
        8'b10111000, // Color (8, 6, 12) (13, 3)
        8'b10110110, // Color (7, 5, 11) (14, 3)
        8'b10110110, // Color (7, 5, 11) (15, 3)
        8'b10110110, // Color (7, 5, 11) (0, 4)
        8'b10111000, // Color (8, 6, 12) (1, 4)
        8'b10111010, // Color (12, 9, 15) (2, 4)
        8'b10110110, // Color (7, 5, 11) (3, 4)
        8'b11000000, // Color (5, 3, 9) (4, 4)
        8'b10110100, // Color (6, 4, 9) (5, 4)
        8'b10110100, // Color (6, 4, 9) (6, 4)
        8'b10110100, // Color (6, 4, 9) (7, 4)
        8'b10110110, // Color (7, 5, 11) (8, 4)
        8'b10111000, // Color (8, 6, 12) (9, 4)
        8'b10110100, // Color (6, 4, 9) (10, 4)
        8'b10110110, // Color (7, 5, 11) (11, 4)
        8'b10111000, // Color (8, 6, 12) (12, 4)
        8'b10110100, // Color (6, 4, 9) (13, 4)
        8'b11000000, // Color (5, 3, 9) (14, 4)
        8'b10110110, // Color (7, 5, 11) (15, 4)
        8'b10111000, // Color (8, 6, 12) (0, 5)
        8'b10111110, // Color (10, 7, 15) (1, 5)
        8'b10111100, // Color (15, 12, 14) (2, 5)
        8'b10111000, // Color (8, 6, 12) (3, 5)
        8'b10110110, // Color (7, 5, 11) (4, 5)
        8'b10110100, // Color (6, 4, 9) (5, 5)
        8'b10110110, // Color (7, 5, 11) (6, 5)
        8'b10110110, // Color (7, 5, 11) (7, 5)
        8'b10111110, // Color (10, 7, 15) (8, 5)
        8'b10111010, // Color (12, 9, 15) (9, 5)
        8'b10111000, // Color (8, 6, 12) (10, 5)
        8'b10110110, // Color (7, 5, 11) (11, 5)
        8'b10110110, // Color (7, 5, 11) (12, 5)
        8'b11000000, // Color (5, 3, 9) (13, 5)
        8'b10110100, // Color (6, 4, 9) (14, 5)
        8'b10110100, // Color (6, 4, 9) (15, 5)
        8'b10111010, // Color (12, 9, 15) (0, 6)
        8'b10111100, // Color (15, 12, 14) (1, 6)
        8'b10111100, // Color (15, 12, 14) (2, 6)
        8'b10111110, // Color (10, 7, 15) (3, 6)
        8'b10111110, // Color (10, 7, 15) (4, 6)
        8'b10110110, // Color (7, 5, 11) (5, 6)
        8'b10110110, // Color (7, 5, 11) (6, 6)
        8'b10110100, // Color (6, 4, 9) (7, 6)
        8'b10110110, // Color (7, 5, 11) (8, 6)
        8'b10111000, // Color (8, 6, 12) (9, 6)
        8'b10110100, // Color (6, 4, 9) (10, 6)
        8'b10110110, // Color (7, 5, 11) (11, 6)
        8'b10110100, // Color (6, 4, 9) (12, 6)
        8'b10110100, // Color (6, 4, 9) (13, 6)
        8'b10110100, // Color (6, 4, 9) (14, 6)
        8'b10111000, // Color (8, 6, 12) (15, 6)
        8'b10110110, // Color (7, 5, 11) (0, 7)
        8'b10111000, // Color (8, 6, 12) (1, 7)
        8'b10111110, // Color (10, 7, 15) (2, 7)
        8'b10110100, // Color (6, 4, 9) (3, 7)
        8'b10110100, // Color (6, 4, 9) (4, 7)
        8'b10110110, // Color (7, 5, 11) (5, 7)
        8'b10111110, // Color (10, 7, 15) (6, 7)
        8'b10110110, // Color (7, 5, 11) (7, 7)
        8'b10111000, // Color (8, 6, 12) (8, 7)
        8'b10110110, // Color (7, 5, 11) (9, 7)
        8'b10110110, // Color (7, 5, 11) (10, 7)
        8'b10111000, // Color (8, 6, 12) (11, 7)
        8'b10110110, // Color (7, 5, 11) (12, 7)
        8'b10110100, // Color (6, 4, 9) (13, 7)
        8'b10111000, // Color (8, 6, 12) (14, 7)
        8'b10110100, // Color (6, 4, 9) (15, 7)
        8'b10110100, // Color (6, 4, 9) (0, 8)
        8'b10110110, // Color (7, 5, 11) (1, 8)
        8'b10111110, // Color (10, 7, 15) (2, 8)
        8'b10110100, // Color (6, 4, 9) (3, 8)
        8'b10111000, // Color (8, 6, 12) (4, 8)
        8'b10111110, // Color (10, 7, 15) (5, 8)
        8'b10111010, // Color (12, 9, 15) (6, 8)
        8'b10111000, // Color (8, 6, 12) (7, 8)
        8'b10110110, // Color (7, 5, 11) (8, 8)
        8'b10110100, // Color (6, 4, 9) (9, 8)
        8'b10110100, // Color (6, 4, 9) (10, 8)
        8'b10110110, // Color (7, 5, 11) (11, 8)
        8'b10110100, // Color (6, 4, 9) (12, 8)
        8'b10111000, // Color (8, 6, 12) (13, 8)
        8'b10111110, // Color (10, 7, 15) (14, 8)
        8'b10110100, // Color (6, 4, 9) (15, 8)
        8'b10110110, // Color (7, 5, 11) (0, 9)
        8'b10110110, // Color (7, 5, 11) (1, 9)
        8'b10110110, // Color (7, 5, 11) (2, 9)
        8'b10111000, // Color (8, 6, 12) (3, 9)
        8'b10111110, // Color (10, 7, 15) (4, 9)
        8'b10110110, // Color (7, 5, 11) (5, 9)
        8'b10111000, // Color (8, 6, 12) (6, 9)
        8'b10110100, // Color (6, 4, 9) (7, 9)
        8'b11000000, // Color (5, 3, 9) (8, 9)
        8'b11000000, // Color (5, 3, 9) (9, 9)
        8'b10110110, // Color (7, 5, 11) (10, 9)
        8'b10111000, // Color (8, 6, 12) (11, 9)
        8'b10110110, // Color (7, 5, 11) (12, 9)
        8'b10111110, // Color (10, 7, 15) (13, 9)
        8'b10111010, // Color (12, 9, 15) (14, 9)
        8'b10111000, // Color (8, 6, 12) (15, 9)
        8'b10110110, // Color (7, 5, 11) (0, 10)
        8'b10110110, // Color (7, 5, 11) (1, 10)
        8'b10111000, // Color (8, 6, 12) (2, 10)
        8'b10111110, // Color (10, 7, 15) (3, 10)
        8'b10111010, // Color (12, 9, 15) (4, 10)
        8'b10111000, // Color (8, 6, 12) (5, 10)
        8'b10110110, // Color (7, 5, 11) (6, 10)
        8'b11000000, // Color (5, 3, 9) (7, 10)
        8'b10110100, // Color (6, 4, 9) (8, 10)
        8'b10110110, // Color (7, 5, 11) (9, 10)
        8'b10111000, // Color (8, 6, 12) (10, 10)
        8'b10111110, // Color (10, 7, 15) (11, 10)
        8'b10111000, // Color (8, 6, 12) (12, 10)
        8'b10110110, // Color (7, 5, 11) (13, 10)
        8'b10111000, // Color (8, 6, 12) (14, 10)
        8'b10110100, // Color (6, 4, 9) (15, 10)
        8'b10110110, // Color (7, 5, 11) (0, 11)
        8'b10111000, // Color (8, 6, 12) (1, 11)
        8'b10111110, // Color (10, 7, 15) (2, 11)
        8'b10111110, // Color (10, 7, 15) (3, 11)
        8'b10111010, // Color (12, 9, 15) (4, 11)
        8'b10111110, // Color (10, 7, 15) (5, 11)
        8'b10111000, // Color (8, 6, 12) (6, 11)
        8'b10110100, // Color (6, 4, 9) (7, 11)
        8'b10110110, // Color (7, 5, 11) (8, 11)
        8'b10111000, // Color (8, 6, 12) (9, 11)
        8'b10111110, // Color (10, 7, 15) (10, 11)
        8'b10111010, // Color (12, 9, 15) (11, 11)
        8'b10111110, // Color (10, 7, 15) (12, 11)
        8'b10111000, // Color (8, 6, 12) (13, 11)
        8'b10110110, // Color (7, 5, 11) (14, 11)
        8'b10110100, // Color (6, 4, 9) (15, 11)
        8'b10110100, // Color (6, 4, 9) (0, 12)
        8'b10111110, // Color (10, 7, 15) (1, 12)
        8'b10111010, // Color (12, 9, 15) (2, 12)
        8'b10111100, // Color (15, 12, 14) (3, 12)
        8'b10111100, // Color (15, 12, 14) (4, 12)
        8'b10111110, // Color (10, 7, 15) (5, 12)
        8'b10111110, // Color (10, 7, 15) (6, 12)
        8'b10110110, // Color (7, 5, 11) (7, 12)
        8'b10110100, // Color (6, 4, 9) (8, 12)
        8'b10110100, // Color (6, 4, 9) (9, 12)
        8'b10110110, // Color (7, 5, 11) (10, 12)
        8'b10111110, // Color (10, 7, 15) (11, 12)
        8'b11000000, // Color (5, 3, 9) (12, 12)
        8'b10110100, // Color (6, 4, 9) (13, 12)
        8'b10111110, // Color (10, 7, 15) (14, 12)
        8'b10110110, // Color (7, 5, 11) (15, 12)
        8'b10110100, // Color (6, 4, 9) (0, 13)
        8'b10110110, // Color (7, 5, 11) (1, 13)
        8'b10111000, // Color (8, 6, 12) (2, 13)
        8'b10111000, // Color (8, 6, 12) (3, 13)
        8'b10111010, // Color (12, 9, 15) (4, 13)
        8'b11000000, // Color (5, 3, 9) (5, 13)
        8'b10110100, // Color (6, 4, 9) (6, 13)
        8'b10110100, // Color (6, 4, 9) (7, 13)
        8'b11000000, // Color (5, 3, 9) (8, 13)
        8'b10110110, // Color (7, 5, 11) (9, 13)
        8'b10110110, // Color (7, 5, 11) (10, 13)
        8'b10110110, // Color (7, 5, 11) (11, 13)
        8'b10110100, // Color (6, 4, 9) (12, 13)
        8'b10110110, // Color (7, 5, 11) (13, 13)
        8'b10111010, // Color (12, 9, 15) (14, 13)
        8'b10111000, // Color (8, 6, 12) (15, 13)
        8'b10110110, // Color (7, 5, 11) (0, 14)
        8'b10110100, // Color (6, 4, 9) (1, 14)
        8'b10110110, // Color (7, 5, 11) (2, 14)
        8'b10111000, // Color (8, 6, 12) (3, 14)
        8'b10111110, // Color (10, 7, 15) (4, 14)
        8'b10110100, // Color (6, 4, 9) (5, 14)
        8'b10110110, // Color (7, 5, 11) (6, 14)
        8'b10110100, // Color (6, 4, 9) (7, 14)
        8'b10110110, // Color (7, 5, 11) (8, 14)
        8'b10111010, // Color (12, 9, 15) (9, 14)
        8'b10110110, // Color (7, 5, 11) (10, 14)
        8'b10110100, // Color (6, 4, 9) (11, 14)
        8'b10110110, // Color (7, 5, 11) (12, 14)
        8'b10111010, // Color (12, 9, 15) (13, 14)
        8'b10111100, // Color (15, 12, 14) (14, 14)
        8'b10111110, // Color (10, 7, 15) (15, 14)
        8'b11000000, // Color (5, 3, 9) (0, 15)
        8'b10110100, // Color (6, 4, 9) (1, 15)
        8'b10110100, // Color (6, 4, 9) (2, 15)
        8'b10110110, // Color (7, 5, 11) (3, 15)
        8'b10111000, // Color (8, 6, 12) (4, 15)
        8'b10110110, // Color (7, 5, 11) (5, 15)
        8'b10110110, // Color (7, 5, 11) (6, 15)
        8'b10110110, // Color (7, 5, 11) (7, 15)
        8'b10111010, // Color (12, 9, 15) (8, 15)
        8'b10111100, // Color (15, 12, 14) (9, 15)
        8'b10111000, // Color (8, 6, 12) (10, 15)
        8'b10110110, // Color (7, 5, 11) (11, 15)
        8'b11000000, // Color (5, 3, 9) (12, 15)
        8'b10110110, // Color (7, 5, 11) (13, 15)
        8'b10111010, // Color (12, 9, 15) (14, 15)
        8'b11000000, // Color (5, 3, 9) (15, 15)
    };

    logic [15:0] texture_address;
    logic [7:0] rom_data;

    always_comb begin
       texture_address = (id << 8) | (y << 4) | x;
    end

    always_ff @(posedge clk) begin
       rom_data <= TEXTURE_ROM[texture_address];
    end

    assign data = rom_data;

endmodule
